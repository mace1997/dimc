// author Mace

module SNAX_DIMC # (
    parameter int unsigned NarrowDataWidth = 64,
    parameter int unsigned WideDataWidth   = 512,
    parameter int unsigned RegAddrWidth    = 32,
    parameter int unsigned RegDataWidth    = 32
)(
    /**************************************************************************/
    // Clock and reset
    /**************************************************************************/
    input  logic                       clk_i,
    input  logic                       rst_ni,

    /**************************************************************************/
    // Accelerator ports
    /**************************************************************************/
    // Ports from accelerator to streamer by writer data movers
    output logic [WideDataWidth-1:0]   acc2stream_0_data_o,
    output logic                       acc2stream_0_valid_o,
    input  logic                       acc2stream_0_ready_i,
    
    // Ports from streamer to accelerator by reader data movers
    input  logic [WideDataWidth-1:0]   stream2acc_0_data_i,
    input  logic                       stream2acc_0_valid_i,
    output logic                       stream2acc_0_ready_o,

    input  logic [WideDataWidth-1:0]   stream2acc_1_data_i,
    input  logic                       stream2acc_1_valid_i,
    output logic                       stream2acc_1_ready_o,

    input  logic [WideDataWidth-1:0]   stream2acc_2_data_i,
    input  logic                       stream2acc_2_valid_i,
    output logic                       stream2acc_2_ready_o,

    input  logic [WideDataWidth-1:0]   stream2acc_3_data_i,
    input  logic                       stream2acc_3_valid_i,
    output logic                       stream2acc_3_ready_o,

    //-----------------------------
    // CSR control ports
    //-----------------------------
    // Request
    input  logic [   RegAddrWidth-1:0] csr_req_addr_i,
    input  logic [   RegDataWidth-1:0] csr_req_data_i,
    input  logic                       csr_req_write_i,
    input  logic                       csr_req_valid_i,
    output logic                       csr_req_ready_o,
    // Response
    output logic [   RegDataWidth-1:0] csr_rsp_data_o,
    output logic                       csr_rsp_valid_o,
    input  logic                       csr_rsp_ready_i
);

// Internal signals

wire rst;

assign rst = ~rst_ni;

wire [11:0] QKV_cal_result_in_0_0, QKV_cal_result_in_0_1, QKV_cal_result_in_0_2, QKV_cal_result_in_0_3, QKV_cal_result_in_0_4, QKV_cal_result_in_0_5, QKV_cal_result_in_0_6, QKV_cal_result_in_0_7, QKV_cal_result_in_0_8, QKV_cal_result_in_0_9, QKV_cal_result_in_0_10, QKV_cal_result_in_0_11, QKV_cal_result_in_0_12, QKV_cal_result_in_0_13, QKV_cal_result_in_0_14, QKV_cal_result_in_0_15,
            QKV_cal_result_in_1_0, QKV_cal_result_in_1_1, QKV_cal_result_in_1_2, QKV_cal_result_in_1_3, QKV_cal_result_in_1_4, QKV_cal_result_in_1_5, QKV_cal_result_in_1_6, QKV_cal_result_in_1_7, QKV_cal_result_in_1_8, QKV_cal_result_in_1_9, QKV_cal_result_in_1_10, QKV_cal_result_in_1_11, QKV_cal_result_in_1_12, QKV_cal_result_in_1_13, QKV_cal_result_in_1_14, QKV_cal_result_in_1_15,
            QKV_cal_result_in_2_0, QKV_cal_result_in_2_1, QKV_cal_result_in_2_2, QKV_cal_result_in_2_3, QKV_cal_result_in_2_4, QKV_cal_result_in_2_5, QKV_cal_result_in_2_6, QKV_cal_result_in_2_7, QKV_cal_result_in_2_8, QKV_cal_result_in_2_9, QKV_cal_result_in_2_10, QKV_cal_result_in_2_11, QKV_cal_result_in_2_12, QKV_cal_result_in_2_13, QKV_cal_result_in_2_14, QKV_cal_result_in_2_15,
            QKV_cal_result_in_3_0, QKV_cal_result_in_3_1, QKV_cal_result_in_3_2, QKV_cal_result_in_3_3, QKV_cal_result_in_3_4, QKV_cal_result_in_3_5, QKV_cal_result_in_3_6, QKV_cal_result_in_3_7, QKV_cal_result_in_3_8, QKV_cal_result_in_3_9, QKV_cal_result_in_3_10, QKV_cal_result_in_3_11, QKV_cal_result_in_3_12, QKV_cal_result_in_3_13, QKV_cal_result_in_3_14, QKV_cal_result_in_3_15,
            QKV_cal_result_in_4_0, QKV_cal_result_in_4_1, QKV_cal_result_in_4_2, QKV_cal_result_in_4_3, QKV_cal_result_in_4_4, QKV_cal_result_in_4_5, QKV_cal_result_in_4_6, QKV_cal_result_in_4_7, QKV_cal_result_in_4_8, QKV_cal_result_in_4_9, QKV_cal_result_in_4_10, QKV_cal_result_in_4_11, QKV_cal_result_in_4_12, QKV_cal_result_in_4_13, QKV_cal_result_in_4_14, QKV_cal_result_in_4_15,
            QKV_cal_result_in_5_0, QKV_cal_result_in_5_1, QKV_cal_result_in_5_2, QKV_cal_result_in_5_3, QKV_cal_result_in_5_4, QKV_cal_result_in_5_5, QKV_cal_result_in_5_6, QKV_cal_result_in_5_7, QKV_cal_result_in_5_8, QKV_cal_result_in_5_9, QKV_cal_result_in_5_10, QKV_cal_result_in_5_11, QKV_cal_result_in_5_12, QKV_cal_result_in_5_13, QKV_cal_result_in_5_14, QKV_cal_result_in_5_15,
            QKV_cal_result_in_6_0, QKV_cal_result_in_6_1, QKV_cal_result_in_6_2, QKV_cal_result_in_6_3, QKV_cal_result_in_6_4, QKV_cal_result_in_6_5, QKV_cal_result_in_6_6, QKV_cal_result_in_6_7, QKV_cal_result_in_6_8, QKV_cal_result_in_6_9, QKV_cal_result_in_6_10, QKV_cal_result_in_6_11, QKV_cal_result_in_6_12, QKV_cal_result_in_6_13, QKV_cal_result_in_6_14, QKV_cal_result_in_6_15,
            QKV_cal_result_in_7_0, QKV_cal_result_in_7_1, QKV_cal_result_in_7_2, QKV_cal_result_in_7_3, QKV_cal_result_in_7_4, QKV_cal_result_in_7_5, QKV_cal_result_in_7_6, QKV_cal_result_in_7_7, QKV_cal_result_in_7_8, QKV_cal_result_in_7_9, QKV_cal_result_in_7_10, QKV_cal_result_in_7_11, QKV_cal_result_in_7_12, QKV_cal_result_in_7_13, QKV_cal_result_in_7_14, QKV_cal_result_in_7_15,
            QKV_cal_result_in_8_0, QKV_cal_result_in_8_1, QKV_cal_result_in_8_2, QKV_cal_result_in_8_3, QKV_cal_result_in_8_4, QKV_cal_result_in_8_5, QKV_cal_result_in_8_6, QKV_cal_result_in_8_7, QKV_cal_result_in_8_8, QKV_cal_result_in_8_9, QKV_cal_result_in_8_10, QKV_cal_result_in_8_11, QKV_cal_result_in_8_12, QKV_cal_result_in_8_13, QKV_cal_result_in_8_14, QKV_cal_result_in_8_15,
            QKV_cal_result_in_9_0, QKV_cal_result_in_9_1, QKV_cal_result_in_9_2, QKV_cal_result_in_9_3, QKV_cal_result_in_9_4, QKV_cal_result_in_9_5, QKV_cal_result_in_9_6, QKV_cal_result_in_9_7, QKV_cal_result_in_9_8, QKV_cal_result_in_9_9, QKV_cal_result_in_9_10, QKV_cal_result_in_9_11, QKV_cal_result_in_9_12, QKV_cal_result_in_9_13, QKV_cal_result_in_9_14, QKV_cal_result_in_9_15,
            QKV_cal_result_in_10_0, QKV_cal_result_in_10_1, QKV_cal_result_in_10_2, QKV_cal_result_in_10_3, QKV_cal_result_in_10_4, QKV_cal_result_in_10_5, QKV_cal_result_in_10_6, QKV_cal_result_in_10_7, QKV_cal_result_in_10_8, QKV_cal_result_in_10_9, QKV_cal_result_in_10_10, QKV_cal_result_in_10_11, QKV_cal_result_in_10_12, QKV_cal_result_in_10_13, QKV_cal_result_in_10_14, QKV_cal_result_in_10_15,
            QKV_cal_result_in_11_0, QKV_cal_result_in_11_1, QKV_cal_result_in_11_2, QKV_cal_result_in_11_3, QKV_cal_result_in_11_4, QKV_cal_result_in_11_5, QKV_cal_result_in_11_6, QKV_cal_result_in_11_7, QKV_cal_result_in_11_8, QKV_cal_result_in_11_9, QKV_cal_result_in_11_10, QKV_cal_result_in_11_11, QKV_cal_result_in_11_12, QKV_cal_result_in_11_13, QKV_cal_result_in_11_14, QKV_cal_result_in_11_15,
            QKV_cal_result_in_12_0, QKV_cal_result_in_12_1, QKV_cal_result_in_12_2, QKV_cal_result_in_12_3, QKV_cal_result_in_12_4, QKV_cal_result_in_12_5, QKV_cal_result_in_12_6, QKV_cal_result_in_12_7, QKV_cal_result_in_12_8, QKV_cal_result_in_12_9, QKV_cal_result_in_12_10, QKV_cal_result_in_12_11, QKV_cal_result_in_12_12, QKV_cal_result_in_12_13, QKV_cal_result_in_12_14, QKV_cal_result_in_12_15,
            QKV_cal_result_in_13_0, QKV_cal_result_in_13_1, QKV_cal_result_in_13_2, QKV_cal_result_in_13_3, QKV_cal_result_in_13_4, QKV_cal_result_in_13_5, QKV_cal_result_in_13_6, QKV_cal_result_in_13_7, QKV_cal_result_in_13_8, QKV_cal_result_in_13_9, QKV_cal_result_in_13_10, QKV_cal_result_in_13_11, QKV_cal_result_in_13_12, QKV_cal_result_in_13_13, QKV_cal_result_in_13_14, QKV_cal_result_in_13_15,
            QKV_cal_result_in_14_0, QKV_cal_result_in_14_1, QKV_cal_result_in_14_2, QKV_cal_result_in_14_3, QKV_cal_result_in_14_4, QKV_cal_result_in_14_5, QKV_cal_result_in_14_6, QKV_cal_result_in_14_7, QKV_cal_result_in_14_8, QKV_cal_result_in_14_9, QKV_cal_result_in_14_10, QKV_cal_result_in_14_11, QKV_cal_result_in_14_12, QKV_cal_result_in_14_13, QKV_cal_result_in_14_14, QKV_cal_result_in_14_15,
            QKV_cal_result_in_15_0, QKV_cal_result_in_15_1, QKV_cal_result_in_15_2, QKV_cal_result_in_15_3, QKV_cal_result_in_15_4, QKV_cal_result_in_15_5, QKV_cal_result_in_15_6, QKV_cal_result_in_15_7, QKV_cal_result_in_15_8, QKV_cal_result_in_15_9, QKV_cal_result_in_15_10, QKV_cal_result_in_15_11, QKV_cal_result_in_15_12, QKV_cal_result_in_15_13, QKV_cal_result_in_15_14, QKV_cal_result_in_15_15,
            QKV_cal_result_in_16_0, QKV_cal_result_in_16_1, QKV_cal_result_in_16_2, QKV_cal_result_in_16_3, QKV_cal_result_in_16_4, QKV_cal_result_in_16_5, QKV_cal_result_in_16_6, QKV_cal_result_in_16_7, QKV_cal_result_in_16_8, QKV_cal_result_in_16_9, QKV_cal_result_in_16_10, QKV_cal_result_in_16_11, QKV_cal_result_in_16_12, QKV_cal_result_in_16_13, QKV_cal_result_in_16_14, QKV_cal_result_in_16_15,
            QKV_cal_result_in_17_0, QKV_cal_result_in_17_1, QKV_cal_result_in_17_2, QKV_cal_result_in_17_3, QKV_cal_result_in_17_4, QKV_cal_result_in_17_5, QKV_cal_result_in_17_6, QKV_cal_result_in_17_7, QKV_cal_result_in_17_8, QKV_cal_result_in_17_9, QKV_cal_result_in_17_10, QKV_cal_result_in_17_11, QKV_cal_result_in_17_12, QKV_cal_result_in_17_13, QKV_cal_result_in_17_14, QKV_cal_result_in_17_15,
            QKV_cal_result_in_18_0, QKV_cal_result_in_18_1, QKV_cal_result_in_18_2, QKV_cal_result_in_18_3, QKV_cal_result_in_18_4, QKV_cal_result_in_18_5, QKV_cal_result_in_18_6, QKV_cal_result_in_18_7, QKV_cal_result_in_18_8, QKV_cal_result_in_18_9, QKV_cal_result_in_18_10, QKV_cal_result_in_18_11, QKV_cal_result_in_18_12, QKV_cal_result_in_18_13, QKV_cal_result_in_18_14, QKV_cal_result_in_18_15,
            QKV_cal_result_in_19_0, QKV_cal_result_in_19_1, QKV_cal_result_in_19_2, QKV_cal_result_in_19_3, QKV_cal_result_in_19_4, QKV_cal_result_in_19_5, QKV_cal_result_in_19_6, QKV_cal_result_in_19_7, QKV_cal_result_in_19_8, QKV_cal_result_in_19_9, QKV_cal_result_in_19_10, QKV_cal_result_in_19_11, QKV_cal_result_in_19_12, QKV_cal_result_in_19_13, QKV_cal_result_in_19_14, QKV_cal_result_in_19_15,
            QKV_cal_result_in_20_0, QKV_cal_result_in_20_1, QKV_cal_result_in_20_2, QKV_cal_result_in_20_3, QKV_cal_result_in_20_4, QKV_cal_result_in_20_5, QKV_cal_result_in_20_6, QKV_cal_result_in_20_7, QKV_cal_result_in_20_8, QKV_cal_result_in_20_9, QKV_cal_result_in_20_10, QKV_cal_result_in_20_11, QKV_cal_result_in_20_12, QKV_cal_result_in_20_13, QKV_cal_result_in_20_14, QKV_cal_result_in_20_15,
            QKV_cal_result_in_21_0, QKV_cal_result_in_21_1, QKV_cal_result_in_21_2, QKV_cal_result_in_21_3, QKV_cal_result_in_21_4, QKV_cal_result_in_21_5, QKV_cal_result_in_21_6, QKV_cal_result_in_21_7, QKV_cal_result_in_21_8, QKV_cal_result_in_21_9, QKV_cal_result_in_21_10, QKV_cal_result_in_21_11, QKV_cal_result_in_21_12, QKV_cal_result_in_21_13, QKV_cal_result_in_21_14, QKV_cal_result_in_21_15,
            QKV_cal_result_in_22_0, QKV_cal_result_in_22_1, QKV_cal_result_in_22_2, QKV_cal_result_in_22_3, QKV_cal_result_in_22_4, QKV_cal_result_in_22_5, QKV_cal_result_in_22_6, QKV_cal_result_in_22_7, QKV_cal_result_in_22_8, QKV_cal_result_in_22_9, QKV_cal_result_in_22_10, QKV_cal_result_in_22_11, QKV_cal_result_in_22_12, QKV_cal_result_in_22_13, QKV_cal_result_in_22_14, QKV_cal_result_in_22_15,
            QKV_cal_result_in_23_0, QKV_cal_result_in_23_1, QKV_cal_result_in_23_2, QKV_cal_result_in_23_3, QKV_cal_result_in_23_4, QKV_cal_result_in_23_5, QKV_cal_result_in_23_6, QKV_cal_result_in_23_7, QKV_cal_result_in_23_8, QKV_cal_result_in_23_9, QKV_cal_result_in_23_10, QKV_cal_result_in_23_11, QKV_cal_result_in_23_12, QKV_cal_result_in_23_13, QKV_cal_result_in_23_14, QKV_cal_result_in_23_15,
            QKV_cal_result_in_24_0, QKV_cal_result_in_24_1, QKV_cal_result_in_24_2, QKV_cal_result_in_24_3, QKV_cal_result_in_24_4, QKV_cal_result_in_24_5, QKV_cal_result_in_24_6, QKV_cal_result_in_24_7, QKV_cal_result_in_24_8, QKV_cal_result_in_24_9, QKV_cal_result_in_24_10, QKV_cal_result_in_24_11, QKV_cal_result_in_24_12, QKV_cal_result_in_24_13, QKV_cal_result_in_24_14, QKV_cal_result_in_24_15,
            QKV_cal_result_in_25_0, QKV_cal_result_in_25_1, QKV_cal_result_in_25_2, QKV_cal_result_in_25_3, QKV_cal_result_in_25_4, QKV_cal_result_in_25_5, QKV_cal_result_in_25_6, QKV_cal_result_in_25_7, QKV_cal_result_in_25_8, QKV_cal_result_in_25_9, QKV_cal_result_in_25_10, QKV_cal_result_in_25_11, QKV_cal_result_in_25_12, QKV_cal_result_in_25_13, QKV_cal_result_in_25_14, QKV_cal_result_in_25_15,
            QKV_cal_result_in_26_0, QKV_cal_result_in_26_1, QKV_cal_result_in_26_2, QKV_cal_result_in_26_3, QKV_cal_result_in_26_4, QKV_cal_result_in_26_5, QKV_cal_result_in_26_6, QKV_cal_result_in_26_7, QKV_cal_result_in_26_8, QKV_cal_result_in_26_9, QKV_cal_result_in_26_10, QKV_cal_result_in_26_11, QKV_cal_result_in_26_12, QKV_cal_result_in_26_13, QKV_cal_result_in_26_14, QKV_cal_result_in_26_15,
            QKV_cal_result_in_27_0, QKV_cal_result_in_27_1, QKV_cal_result_in_27_2, QKV_cal_result_in_27_3, QKV_cal_result_in_27_4, QKV_cal_result_in_27_5, QKV_cal_result_in_27_6, QKV_cal_result_in_27_7, QKV_cal_result_in_27_8, QKV_cal_result_in_27_9, QKV_cal_result_in_27_10, QKV_cal_result_in_27_11, QKV_cal_result_in_27_12, QKV_cal_result_in_27_13, QKV_cal_result_in_27_14, QKV_cal_result_in_27_15,
            QKV_cal_result_in_28_0, QKV_cal_result_in_28_1, QKV_cal_result_in_28_2, QKV_cal_result_in_28_3, QKV_cal_result_in_28_4, QKV_cal_result_in_28_5, QKV_cal_result_in_28_6, QKV_cal_result_in_28_7, QKV_cal_result_in_28_8, QKV_cal_result_in_28_9, QKV_cal_result_in_28_10, QKV_cal_result_in_28_11, QKV_cal_result_in_28_12, QKV_cal_result_in_28_13, QKV_cal_result_in_28_14, QKV_cal_result_in_28_15,
            QKV_cal_result_in_29_0, QKV_cal_result_in_29_1, QKV_cal_result_in_29_2, QKV_cal_result_in_29_3, QKV_cal_result_in_29_4, QKV_cal_result_in_29_5, QKV_cal_result_in_29_6, QKV_cal_result_in_29_7, QKV_cal_result_in_29_8, QKV_cal_result_in_29_9, QKV_cal_result_in_29_10, QKV_cal_result_in_29_11, QKV_cal_result_in_29_12, QKV_cal_result_in_29_13, QKV_cal_result_in_29_14, QKV_cal_result_in_29_15,
            QKV_cal_result_in_30_0, QKV_cal_result_in_30_1, QKV_cal_result_in_30_2, QKV_cal_result_in_30_3, QKV_cal_result_in_30_4, QKV_cal_result_in_30_5, QKV_cal_result_in_30_6, QKV_cal_result_in_30_7, QKV_cal_result_in_30_8, QKV_cal_result_in_30_9, QKV_cal_result_in_30_10, QKV_cal_result_in_30_11, QKV_cal_result_in_30_12, QKV_cal_result_in_30_13, QKV_cal_result_in_30_14, QKV_cal_result_in_30_15,
            QKV_cal_result_in_31_0, QKV_cal_result_in_31_1, QKV_cal_result_in_31_2, QKV_cal_result_in_31_3, QKV_cal_result_in_31_4, QKV_cal_result_in_31_5, QKV_cal_result_in_31_6, QKV_cal_result_in_31_7, QKV_cal_result_in_31_8, QKV_cal_result_in_31_9, QKV_cal_result_in_31_10, QKV_cal_result_in_31_11, QKV_cal_result_in_31_12, QKV_cal_result_in_31_13, QKV_cal_result_in_31_14, QKV_cal_result_in_31_15;

wire [11:0] QKT_cal_result_in_0_0, QKT_cal_result_in_0_1, QKT_cal_result_in_0_2, QKT_cal_result_in_0_3, QKT_cal_result_in_0_4, QKT_cal_result_in_0_5, QKT_cal_result_in_0_6, QKT_cal_result_in_0_7, QKT_cal_result_in_0_8, QKT_cal_result_in_0_9, QKT_cal_result_in_0_10, QKT_cal_result_in_0_11, QKT_cal_result_in_0_12, QKT_cal_result_in_0_13, QKT_cal_result_in_0_14, QKT_cal_result_in_0_15,
            QKT_cal_result_in_1_0, QKT_cal_result_in_1_1, QKT_cal_result_in_1_2, QKT_cal_result_in_1_3, QKT_cal_result_in_1_4, QKT_cal_result_in_1_5, QKT_cal_result_in_1_6, QKT_cal_result_in_1_7, QKT_cal_result_in_1_8, QKT_cal_result_in_1_9, QKT_cal_result_in_1_10, QKT_cal_result_in_1_11, QKT_cal_result_in_1_12, QKT_cal_result_in_1_13, QKT_cal_result_in_1_14, QKT_cal_result_in_1_15,
            QKT_cal_result_in_2_0, QKT_cal_result_in_2_1, QKT_cal_result_in_2_2, QKT_cal_result_in_2_3, QKT_cal_result_in_2_4, QKT_cal_result_in_2_5, QKT_cal_result_in_2_6, QKT_cal_result_in_2_7, QKT_cal_result_in_2_8, QKT_cal_result_in_2_9, QKT_cal_result_in_2_10, QKT_cal_result_in_2_11, QKT_cal_result_in_2_12, QKT_cal_result_in_2_13, QKT_cal_result_in_2_14, QKT_cal_result_in_2_15,
            QKT_cal_result_in_3_0, QKT_cal_result_in_3_1, QKT_cal_result_in_3_2, QKT_cal_result_in_3_3, QKT_cal_result_in_3_4, QKT_cal_result_in_3_5, QKT_cal_result_in_3_6, QKT_cal_result_in_3_7, QKT_cal_result_in_3_8, QKT_cal_result_in_3_9, QKT_cal_result_in_3_10, QKT_cal_result_in_3_11, QKT_cal_result_in_3_12, QKT_cal_result_in_3_13, QKT_cal_result_in_3_14, QKT_cal_result_in_3_15;

wire [5:0] QKV_addr_out_0,  QKV_addr_out_1,  QKV_addr_out_2,  QKV_addr_out_3,  QKV_addr_out_4,  QKV_addr_out_5,  QKV_addr_out_6,  QKV_addr_out_7, 
           QKV_addr_out_8,  QKV_addr_out_9,  QKV_addr_out_10, QKV_addr_out_11, QKV_addr_out_12, QKV_addr_out_13, QKV_addr_out_14, QKV_addr_out_15,
           QKV_addr_out_16, QKV_addr_out_17, QKV_addr_out_18, QKV_addr_out_19, QKV_addr_out_20, QKV_addr_out_21, QKV_addr_out_22, QKV_addr_out_23,
           QKV_addr_out_24, QKV_addr_out_25, QKV_addr_out_26, QKV_addr_out_27, QKV_addr_out_28, QKV_addr_out_29, QKV_addr_out_30, QKV_addr_out_31;

wire [5:0] QKT_addr_out_0, QKT_addr_out_1, QKT_addr_out_2, QKT_addr_out_3;

wire [7:0] QKV_weight_out_0_0, QKV_weight_out_0_1, QKV_weight_out_0_2, QKV_weight_out_0_3, QKV_weight_out_0_4, QKV_weight_out_0_5, QKV_weight_out_0_6, QKV_weight_out_0_7, QKV_weight_out_0_8, QKV_weight_out_0_9, QKV_weight_out_0_10, QKV_weight_out_0_11, QKV_weight_out_0_12, QKV_weight_out_0_13, QKV_weight_out_0_14, QKV_weight_out_0_15, 
           QKV_weight_out_1_0, QKV_weight_out_1_1, QKV_weight_out_1_2, QKV_weight_out_1_3, QKV_weight_out_1_4, QKV_weight_out_1_5, QKV_weight_out_1_6, QKV_weight_out_1_7, QKV_weight_out_1_8, QKV_weight_out_1_9, QKV_weight_out_1_10, QKV_weight_out_1_11, QKV_weight_out_1_12, QKV_weight_out_1_13, QKV_weight_out_1_14, QKV_weight_out_1_15, 
           QKV_weight_out_2_0, QKV_weight_out_2_1, QKV_weight_out_2_2, QKV_weight_out_2_3, QKV_weight_out_2_4, QKV_weight_out_2_5, QKV_weight_out_2_6, QKV_weight_out_2_7, QKV_weight_out_2_8, QKV_weight_out_2_9, QKV_weight_out_2_10, QKV_weight_out_2_11, QKV_weight_out_2_12, QKV_weight_out_2_13, QKV_weight_out_2_14, QKV_weight_out_2_15, 
           QKV_weight_out_3_0, QKV_weight_out_3_1, QKV_weight_out_3_2, QKV_weight_out_3_3, QKV_weight_out_3_4, QKV_weight_out_3_5, QKV_weight_out_3_6, QKV_weight_out_3_7, QKV_weight_out_3_8, QKV_weight_out_3_9, QKV_weight_out_3_10, QKV_weight_out_3_11, QKV_weight_out_3_12, QKV_weight_out_3_13, QKV_weight_out_3_14, QKV_weight_out_3_15, 
           QKV_weight_out_4_0, QKV_weight_out_4_1, QKV_weight_out_4_2, QKV_weight_out_4_3, QKV_weight_out_4_4, QKV_weight_out_4_5, QKV_weight_out_4_6, QKV_weight_out_4_7, QKV_weight_out_4_8, QKV_weight_out_4_9, QKV_weight_out_4_10, QKV_weight_out_4_11, QKV_weight_out_4_12, QKV_weight_out_4_13, QKV_weight_out_4_14, QKV_weight_out_4_15, 
           QKV_weight_out_5_0, QKV_weight_out_5_1, QKV_weight_out_5_2, QKV_weight_out_5_3, QKV_weight_out_5_4, QKV_weight_out_5_5, QKV_weight_out_5_6, QKV_weight_out_5_7, QKV_weight_out_5_8, QKV_weight_out_5_9, QKV_weight_out_5_10, QKV_weight_out_5_11, QKV_weight_out_5_12, QKV_weight_out_5_13, QKV_weight_out_5_14, QKV_weight_out_5_15, 
           QKV_weight_out_6_0, QKV_weight_out_6_1, QKV_weight_out_6_2, QKV_weight_out_6_3, QKV_weight_out_6_4, QKV_weight_out_6_5, QKV_weight_out_6_6, QKV_weight_out_6_7, QKV_weight_out_6_8, QKV_weight_out_6_9, QKV_weight_out_6_10, QKV_weight_out_6_11, QKV_weight_out_6_12, QKV_weight_out_6_13, QKV_weight_out_6_14, QKV_weight_out_6_15, 
           QKV_weight_out_7_0, QKV_weight_out_7_1, QKV_weight_out_7_2, QKV_weight_out_7_3, QKV_weight_out_7_4, QKV_weight_out_7_5, QKV_weight_out_7_6, QKV_weight_out_7_7, QKV_weight_out_7_8, QKV_weight_out_7_9, QKV_weight_out_7_10, QKV_weight_out_7_11, QKV_weight_out_7_12, QKV_weight_out_7_13, QKV_weight_out_7_14, QKV_weight_out_7_15, 
           QKV_weight_out_8_0, QKV_weight_out_8_1, QKV_weight_out_8_2, QKV_weight_out_8_3, QKV_weight_out_8_4, QKV_weight_out_8_5, QKV_weight_out_8_6, QKV_weight_out_8_7, QKV_weight_out_8_8, QKV_weight_out_8_9, QKV_weight_out_8_10, QKV_weight_out_8_11, QKV_weight_out_8_12, QKV_weight_out_8_13, QKV_weight_out_8_14, QKV_weight_out_8_15, 
           QKV_weight_out_9_0, QKV_weight_out_9_1, QKV_weight_out_9_2, QKV_weight_out_9_3, QKV_weight_out_9_4, QKV_weight_out_9_5, QKV_weight_out_9_6, QKV_weight_out_9_7, QKV_weight_out_9_8, QKV_weight_out_9_9, QKV_weight_out_9_10, QKV_weight_out_9_11, QKV_weight_out_9_12, QKV_weight_out_9_13, QKV_weight_out_9_14, QKV_weight_out_9_15, 
           QKV_weight_out_10_0, QKV_weight_out_10_1, QKV_weight_out_10_2, QKV_weight_out_10_3, QKV_weight_out_10_4, QKV_weight_out_10_5, QKV_weight_out_10_6, QKV_weight_out_10_7, QKV_weight_out_10_8, QKV_weight_out_10_9, QKV_weight_out_10_10, QKV_weight_out_10_11, QKV_weight_out_10_12, QKV_weight_out_10_13, QKV_weight_out_10_14, QKV_weight_out_10_15, 
           QKV_weight_out_11_0, QKV_weight_out_11_1, QKV_weight_out_11_2, QKV_weight_out_11_3, QKV_weight_out_11_4, QKV_weight_out_11_5, QKV_weight_out_11_6, QKV_weight_out_11_7, QKV_weight_out_11_8, QKV_weight_out_11_9, QKV_weight_out_11_10, QKV_weight_out_11_11, QKV_weight_out_11_12, QKV_weight_out_11_13, QKV_weight_out_11_14, QKV_weight_out_11_15, 
           QKV_weight_out_12_0, QKV_weight_out_12_1, QKV_weight_out_12_2, QKV_weight_out_12_3, QKV_weight_out_12_4, QKV_weight_out_12_5, QKV_weight_out_12_6, QKV_weight_out_12_7, QKV_weight_out_12_8, QKV_weight_out_12_9, QKV_weight_out_12_10, QKV_weight_out_12_11, QKV_weight_out_12_12, QKV_weight_out_12_13, QKV_weight_out_12_14, QKV_weight_out_12_15, 
           QKV_weight_out_13_0, QKV_weight_out_13_1, QKV_weight_out_13_2, QKV_weight_out_13_3, QKV_weight_out_13_4, QKV_weight_out_13_5, QKV_weight_out_13_6, QKV_weight_out_13_7, QKV_weight_out_13_8, QKV_weight_out_13_9, QKV_weight_out_13_10, QKV_weight_out_13_11, QKV_weight_out_13_12, QKV_weight_out_13_13, QKV_weight_out_13_14, QKV_weight_out_13_15, 
           QKV_weight_out_14_0, QKV_weight_out_14_1, QKV_weight_out_14_2, QKV_weight_out_14_3, QKV_weight_out_14_4, QKV_weight_out_14_5, QKV_weight_out_14_6, QKV_weight_out_14_7, QKV_weight_out_14_8, QKV_weight_out_14_9, QKV_weight_out_14_10, QKV_weight_out_14_11, QKV_weight_out_14_12, QKV_weight_out_14_13, QKV_weight_out_14_14, QKV_weight_out_14_15, 
           QKV_weight_out_15_0, QKV_weight_out_15_1, QKV_weight_out_15_2, QKV_weight_out_15_3, QKV_weight_out_15_4, QKV_weight_out_15_5, QKV_weight_out_15_6, QKV_weight_out_15_7, QKV_weight_out_15_8, QKV_weight_out_15_9, QKV_weight_out_15_10, QKV_weight_out_15_11, QKV_weight_out_15_12, QKV_weight_out_15_13, QKV_weight_out_15_14, QKV_weight_out_15_15, 
           QKV_weight_out_16_0, QKV_weight_out_16_1, QKV_weight_out_16_2, QKV_weight_out_16_3, QKV_weight_out_16_4, QKV_weight_out_16_5, QKV_weight_out_16_6, QKV_weight_out_16_7, QKV_weight_out_16_8, QKV_weight_out_16_9, QKV_weight_out_16_10, QKV_weight_out_16_11, QKV_weight_out_16_12, QKV_weight_out_16_13, QKV_weight_out_16_14, QKV_weight_out_16_15, 
           QKV_weight_out_17_0, QKV_weight_out_17_1, QKV_weight_out_17_2, QKV_weight_out_17_3, QKV_weight_out_17_4, QKV_weight_out_17_5, QKV_weight_out_17_6, QKV_weight_out_17_7, QKV_weight_out_17_8, QKV_weight_out_17_9, QKV_weight_out_17_10, QKV_weight_out_17_11, QKV_weight_out_17_12, QKV_weight_out_17_13, QKV_weight_out_17_14, QKV_weight_out_17_15, 
           QKV_weight_out_18_0, QKV_weight_out_18_1, QKV_weight_out_18_2, QKV_weight_out_18_3, QKV_weight_out_18_4, QKV_weight_out_18_5, QKV_weight_out_18_6, QKV_weight_out_18_7, QKV_weight_out_18_8, QKV_weight_out_18_9, QKV_weight_out_18_10, QKV_weight_out_18_11, QKV_weight_out_18_12, QKV_weight_out_18_13, QKV_weight_out_18_14, QKV_weight_out_18_15, 
           QKV_weight_out_19_0, QKV_weight_out_19_1, QKV_weight_out_19_2, QKV_weight_out_19_3, QKV_weight_out_19_4, QKV_weight_out_19_5, QKV_weight_out_19_6, QKV_weight_out_19_7, QKV_weight_out_19_8, QKV_weight_out_19_9, QKV_weight_out_19_10, QKV_weight_out_19_11, QKV_weight_out_19_12, QKV_weight_out_19_13, QKV_weight_out_19_14, QKV_weight_out_19_15, 
           QKV_weight_out_20_0, QKV_weight_out_20_1, QKV_weight_out_20_2, QKV_weight_out_20_3, QKV_weight_out_20_4, QKV_weight_out_20_5, QKV_weight_out_20_6, QKV_weight_out_20_7, QKV_weight_out_20_8, QKV_weight_out_20_9, QKV_weight_out_20_10, QKV_weight_out_20_11, QKV_weight_out_20_12, QKV_weight_out_20_13, QKV_weight_out_20_14, QKV_weight_out_20_15, 
           QKV_weight_out_21_0, QKV_weight_out_21_1, QKV_weight_out_21_2, QKV_weight_out_21_3, QKV_weight_out_21_4, QKV_weight_out_21_5, QKV_weight_out_21_6, QKV_weight_out_21_7, QKV_weight_out_21_8, QKV_weight_out_21_9, QKV_weight_out_21_10, QKV_weight_out_21_11, QKV_weight_out_21_12, QKV_weight_out_21_13, QKV_weight_out_21_14, QKV_weight_out_21_15, 
           QKV_weight_out_22_0, QKV_weight_out_22_1, QKV_weight_out_22_2, QKV_weight_out_22_3, QKV_weight_out_22_4, QKV_weight_out_22_5, QKV_weight_out_22_6, QKV_weight_out_22_7, QKV_weight_out_22_8, QKV_weight_out_22_9, QKV_weight_out_22_10, QKV_weight_out_22_11, QKV_weight_out_22_12, QKV_weight_out_22_13, QKV_weight_out_22_14, QKV_weight_out_22_15, 
           QKV_weight_out_23_0, QKV_weight_out_23_1, QKV_weight_out_23_2, QKV_weight_out_23_3, QKV_weight_out_23_4, QKV_weight_out_23_5, QKV_weight_out_23_6, QKV_weight_out_23_7, QKV_weight_out_23_8, QKV_weight_out_23_9, QKV_weight_out_23_10, QKV_weight_out_23_11, QKV_weight_out_23_12, QKV_weight_out_23_13, QKV_weight_out_23_14, QKV_weight_out_23_15, 
           QKV_weight_out_24_0, QKV_weight_out_24_1, QKV_weight_out_24_2, QKV_weight_out_24_3, QKV_weight_out_24_4, QKV_weight_out_24_5, QKV_weight_out_24_6, QKV_weight_out_24_7, QKV_weight_out_24_8, QKV_weight_out_24_9, QKV_weight_out_24_10, QKV_weight_out_24_11, QKV_weight_out_24_12, QKV_weight_out_24_13, QKV_weight_out_24_14, QKV_weight_out_24_15, 
           QKV_weight_out_25_0, QKV_weight_out_25_1, QKV_weight_out_25_2, QKV_weight_out_25_3, QKV_weight_out_25_4, QKV_weight_out_25_5, QKV_weight_out_25_6, QKV_weight_out_25_7, QKV_weight_out_25_8, QKV_weight_out_25_9, QKV_weight_out_25_10, QKV_weight_out_25_11, QKV_weight_out_25_12, QKV_weight_out_25_13, QKV_weight_out_25_14, QKV_weight_out_25_15, 
           QKV_weight_out_26_0, QKV_weight_out_26_1, QKV_weight_out_26_2, QKV_weight_out_26_3, QKV_weight_out_26_4, QKV_weight_out_26_5, QKV_weight_out_26_6, QKV_weight_out_26_7, QKV_weight_out_26_8, QKV_weight_out_26_9, QKV_weight_out_26_10, QKV_weight_out_26_11, QKV_weight_out_26_12, QKV_weight_out_26_13, QKV_weight_out_26_14, QKV_weight_out_26_15, 
           QKV_weight_out_27_0, QKV_weight_out_27_1, QKV_weight_out_27_2, QKV_weight_out_27_3, QKV_weight_out_27_4, QKV_weight_out_27_5, QKV_weight_out_27_6, QKV_weight_out_27_7, QKV_weight_out_27_8, QKV_weight_out_27_9, QKV_weight_out_27_10, QKV_weight_out_27_11, QKV_weight_out_27_12, QKV_weight_out_27_13, QKV_weight_out_27_14, QKV_weight_out_27_15, 
           QKV_weight_out_28_0, QKV_weight_out_28_1, QKV_weight_out_28_2, QKV_weight_out_28_3, QKV_weight_out_28_4, QKV_weight_out_28_5, QKV_weight_out_28_6, QKV_weight_out_28_7, QKV_weight_out_28_8, QKV_weight_out_28_9, QKV_weight_out_28_10, QKV_weight_out_28_11, QKV_weight_out_28_12, QKV_weight_out_28_13, QKV_weight_out_28_14, QKV_weight_out_28_15, 
           QKV_weight_out_29_0, QKV_weight_out_29_1, QKV_weight_out_29_2, QKV_weight_out_29_3, QKV_weight_out_29_4, QKV_weight_out_29_5, QKV_weight_out_29_6, QKV_weight_out_29_7, QKV_weight_out_29_8, QKV_weight_out_29_9, QKV_weight_out_29_10, QKV_weight_out_29_11, QKV_weight_out_29_12, QKV_weight_out_29_13, QKV_weight_out_29_14, QKV_weight_out_29_15, 
           QKV_weight_out_30_0, QKV_weight_out_30_1, QKV_weight_out_30_2, QKV_weight_out_30_3, QKV_weight_out_30_4, QKV_weight_out_30_5, QKV_weight_out_30_6, QKV_weight_out_30_7, QKV_weight_out_30_8, QKV_weight_out_30_9, QKV_weight_out_30_10, QKV_weight_out_30_11, QKV_weight_out_30_12, QKV_weight_out_30_13, QKV_weight_out_30_14, QKV_weight_out_30_15, 
           QKV_weight_out_31_0, QKV_weight_out_31_1, QKV_weight_out_31_2, QKV_weight_out_31_3, QKV_weight_out_31_4, QKV_weight_out_31_5, QKV_weight_out_31_6, QKV_weight_out_31_7, QKV_weight_out_31_8, QKV_weight_out_31_9, QKV_weight_out_31_10, QKV_weight_out_31_11, QKV_weight_out_31_12, QKV_weight_out_31_13, QKV_weight_out_31_14, QKV_weight_out_31_15;

wire [7:0] QKT_weight_out_0_0, QKT_weight_out_0_1, QKT_weight_out_0_2, QKT_weight_out_0_3, QKT_weight_out_0_4, QKT_weight_out_0_5, QKT_weight_out_0_6, QKT_weight_out_0_7, QKT_weight_out_0_8, QKT_weight_out_0_9, QKT_weight_out_0_10, QKT_weight_out_0_11, QKT_weight_out_0_12, QKT_weight_out_0_13, QKT_weight_out_0_14, QKT_weight_out_0_15,
           QKT_weight_out_1_0, QKT_weight_out_1_1, QKT_weight_out_1_2, QKT_weight_out_1_3, QKT_weight_out_1_4, QKT_weight_out_1_5, QKT_weight_out_1_6, QKT_weight_out_1_7, QKT_weight_out_1_8, QKT_weight_out_1_9, QKT_weight_out_1_10, QKT_weight_out_1_11, QKT_weight_out_1_12, QKT_weight_out_1_13, QKT_weight_out_1_14, QKT_weight_out_1_15,
           QKT_weight_out_2_0, QKT_weight_out_2_1, QKT_weight_out_2_2, QKT_weight_out_2_3, QKT_weight_out_2_4, QKT_weight_out_2_5, QKT_weight_out_2_6, QKT_weight_out_2_7, QKT_weight_out_2_8, QKT_weight_out_2_9, QKT_weight_out_2_10, QKT_weight_out_2_11, QKT_weight_out_2_12, QKT_weight_out_2_13, QKT_weight_out_2_14, QKT_weight_out_2_15,
           QKT_weight_out_3_0, QKT_weight_out_3_1, QKT_weight_out_3_2, QKT_weight_out_3_3, QKT_weight_out_3_4, QKT_weight_out_3_5, QKT_weight_out_3_6, QKT_weight_out_3_7, QKT_weight_out_3_8, QKT_weight_out_3_9, QKT_weight_out_3_10, QKT_weight_out_3_11, QKT_weight_out_3_12, QKT_weight_out_3_13, QKT_weight_out_3_14, QKT_weight_out_3_15;

wire [3:0] QKV_data_out_0_0, QKV_data_out_0_1, QKV_data_out_0_2, QKV_data_out_0_3, QKV_data_out_0_4, QKV_data_out_0_5, QKV_data_out_0_6, QKV_data_out_0_7, QKV_data_out_0_8, QKV_data_out_0_9, QKV_data_out_0_10, QKV_data_out_0_11, QKV_data_out_0_12, QKV_data_out_0_13, QKV_data_out_0_14, QKV_data_out_0_15,
           QKV_data_out_1_0, QKV_data_out_1_1, QKV_data_out_1_2, QKV_data_out_1_3, QKV_data_out_1_4, QKV_data_out_1_5, QKV_data_out_1_6, QKV_data_out_1_7, QKV_data_out_1_8, QKV_data_out_1_9, QKV_data_out_1_10, QKV_data_out_1_11, QKV_data_out_1_12, QKV_data_out_1_13, QKV_data_out_1_14, QKV_data_out_1_15,
           QKV_data_out_2_0, QKV_data_out_2_1, QKV_data_out_2_2, QKV_data_out_2_3, QKV_data_out_2_4, QKV_data_out_2_5, QKV_data_out_2_6, QKV_data_out_2_7, QKV_data_out_2_8, QKV_data_out_2_9, QKV_data_out_2_10, QKV_data_out_2_11, QKV_data_out_2_12, QKV_data_out_2_13, QKV_data_out_2_14, QKV_data_out_2_15,
           QKV_data_out_3_0, QKV_data_out_3_1, QKV_data_out_3_2, QKV_data_out_3_3, QKV_data_out_3_4, QKV_data_out_3_5, QKV_data_out_3_6, QKV_data_out_3_7, QKV_data_out_3_8, QKV_data_out_3_9, QKV_data_out_3_10, QKV_data_out_3_11, QKV_data_out_3_12, QKV_data_out_3_13, QKV_data_out_3_14, QKV_data_out_3_15,
           QKV_data_out_4_0, QKV_data_out_4_1, QKV_data_out_4_2, QKV_data_out_4_3, QKV_data_out_4_4, QKV_data_out_4_5, QKV_data_out_4_6, QKV_data_out_4_7, QKV_data_out_4_8, QKV_data_out_4_9, QKV_data_out_4_10, QKV_data_out_4_11, QKV_data_out_4_12, QKV_data_out_4_13, QKV_data_out_4_14, QKV_data_out_4_15,
           QKV_data_out_5_0, QKV_data_out_5_1, QKV_data_out_5_2, QKV_data_out_5_3, QKV_data_out_5_4, QKV_data_out_5_5, QKV_data_out_5_6, QKV_data_out_5_7, QKV_data_out_5_8, QKV_data_out_5_9, QKV_data_out_5_10, QKV_data_out_5_11, QKV_data_out_5_12, QKV_data_out_5_13, QKV_data_out_5_14, QKV_data_out_5_15,
           QKV_data_out_6_0, QKV_data_out_6_1, QKV_data_out_6_2, QKV_data_out_6_3, QKV_data_out_6_4, QKV_data_out_6_5, QKV_data_out_6_6, QKV_data_out_6_7, QKV_data_out_6_8, QKV_data_out_6_9, QKV_data_out_6_10, QKV_data_out_6_11, QKV_data_out_6_12, QKV_data_out_6_13, QKV_data_out_6_14, QKV_data_out_6_15,
           QKV_data_out_7_0, QKV_data_out_7_1, QKV_data_out_7_2, QKV_data_out_7_3, QKV_data_out_7_4, QKV_data_out_7_5, QKV_data_out_7_6, QKV_data_out_7_7, QKV_data_out_7_8, QKV_data_out_7_9, QKV_data_out_7_10, QKV_data_out_7_11, QKV_data_out_7_12, QKV_data_out_7_13, QKV_data_out_7_14, QKV_data_out_7_15,
           QKV_data_out_8_0, QKV_data_out_8_1, QKV_data_out_8_2, QKV_data_out_8_3, QKV_data_out_8_4, QKV_data_out_8_5, QKV_data_out_8_6, QKV_data_out_8_7, QKV_data_out_8_8, QKV_data_out_8_9, QKV_data_out_8_10, QKV_data_out_8_11, QKV_data_out_8_12, QKV_data_out_8_13, QKV_data_out_8_14, QKV_data_out_8_15,
           QKV_data_out_9_0, QKV_data_out_9_1, QKV_data_out_9_2, QKV_data_out_9_3, QKV_data_out_9_4, QKV_data_out_9_5, QKV_data_out_9_6, QKV_data_out_9_7, QKV_data_out_9_8, QKV_data_out_9_9, QKV_data_out_9_10, QKV_data_out_9_11, QKV_data_out_9_12, QKV_data_out_9_13, QKV_data_out_9_14, QKV_data_out_9_15,
           QKV_data_out_10_0, QKV_data_out_10_1, QKV_data_out_10_2, QKV_data_out_10_3, QKV_data_out_10_4, QKV_data_out_10_5, QKV_data_out_10_6, QKV_data_out_10_7, QKV_data_out_10_8, QKV_data_out_10_9, QKV_data_out_10_10, QKV_data_out_10_11, QKV_data_out_10_12, QKV_data_out_10_13, QKV_data_out_10_14, QKV_data_out_10_15,
           QKV_data_out_11_0, QKV_data_out_11_1, QKV_data_out_11_2, QKV_data_out_11_3, QKV_data_out_11_4, QKV_data_out_11_5, QKV_data_out_11_6, QKV_data_out_11_7, QKV_data_out_11_8, QKV_data_out_11_9, QKV_data_out_11_10, QKV_data_out_11_11, QKV_data_out_11_12, QKV_data_out_11_13, QKV_data_out_11_14, QKV_data_out_11_15,
           QKV_data_out_12_0, QKV_data_out_12_1, QKV_data_out_12_2, QKV_data_out_12_3, QKV_data_out_12_4, QKV_data_out_12_5, QKV_data_out_12_6, QKV_data_out_12_7, QKV_data_out_12_8, QKV_data_out_12_9, QKV_data_out_12_10, QKV_data_out_12_11, QKV_data_out_12_12, QKV_data_out_12_13, QKV_data_out_12_14, QKV_data_out_12_15,
           QKV_data_out_13_0, QKV_data_out_13_1, QKV_data_out_13_2, QKV_data_out_13_3, QKV_data_out_13_4, QKV_data_out_13_5, QKV_data_out_13_6, QKV_data_out_13_7, QKV_data_out_13_8, QKV_data_out_13_9, QKV_data_out_13_10, QKV_data_out_13_11, QKV_data_out_13_12, QKV_data_out_13_13, QKV_data_out_13_14, QKV_data_out_13_15,
           QKV_data_out_14_0, QKV_data_out_14_1, QKV_data_out_14_2, QKV_data_out_14_3, QKV_data_out_14_4, QKV_data_out_14_5, QKV_data_out_14_6, QKV_data_out_14_7, QKV_data_out_14_8, QKV_data_out_14_9, QKV_data_out_14_10, QKV_data_out_14_11, QKV_data_out_14_12, QKV_data_out_14_13, QKV_data_out_14_14, QKV_data_out_14_15,
           QKV_data_out_15_0, QKV_data_out_15_1, QKV_data_out_15_2, QKV_data_out_15_3, QKV_data_out_15_4, QKV_data_out_15_5, QKV_data_out_15_6, QKV_data_out_15_7, QKV_data_out_15_8, QKV_data_out_15_9, QKV_data_out_15_10, QKV_data_out_15_11, QKV_data_out_15_12, QKV_data_out_15_13, QKV_data_out_15_14, QKV_data_out_15_15,
           QKV_data_out_16_0, QKV_data_out_16_1, QKV_data_out_16_2, QKV_data_out_16_3, QKV_data_out_16_4, QKV_data_out_16_5, QKV_data_out_16_6, QKV_data_out_16_7, QKV_data_out_16_8, QKV_data_out_16_9, QKV_data_out_16_10, QKV_data_out_16_11, QKV_data_out_16_12, QKV_data_out_16_13, QKV_data_out_16_14, QKV_data_out_16_15,
           QKV_data_out_17_0, QKV_data_out_17_1, QKV_data_out_17_2, QKV_data_out_17_3, QKV_data_out_17_4, QKV_data_out_17_5, QKV_data_out_17_6, QKV_data_out_17_7, QKV_data_out_17_8, QKV_data_out_17_9, QKV_data_out_17_10, QKV_data_out_17_11, QKV_data_out_17_12, QKV_data_out_17_13, QKV_data_out_17_14, QKV_data_out_17_15,
           QKV_data_out_18_0, QKV_data_out_18_1, QKV_data_out_18_2, QKV_data_out_18_3, QKV_data_out_18_4, QKV_data_out_18_5, QKV_data_out_18_6, QKV_data_out_18_7, QKV_data_out_18_8, QKV_data_out_18_9, QKV_data_out_18_10, QKV_data_out_18_11, QKV_data_out_18_12, QKV_data_out_18_13, QKV_data_out_18_14, QKV_data_out_18_15,
           QKV_data_out_19_0, QKV_data_out_19_1, QKV_data_out_19_2, QKV_data_out_19_3, QKV_data_out_19_4, QKV_data_out_19_5, QKV_data_out_19_6, QKV_data_out_19_7, QKV_data_out_19_8, QKV_data_out_19_9, QKV_data_out_19_10, QKV_data_out_19_11, QKV_data_out_19_12, QKV_data_out_19_13, QKV_data_out_19_14, QKV_data_out_19_15,
           QKV_data_out_20_0, QKV_data_out_20_1, QKV_data_out_20_2, QKV_data_out_20_3, QKV_data_out_20_4, QKV_data_out_20_5, QKV_data_out_20_6, QKV_data_out_20_7, QKV_data_out_20_8, QKV_data_out_20_9, QKV_data_out_20_10, QKV_data_out_20_11, QKV_data_out_20_12, QKV_data_out_20_13, QKV_data_out_20_14, QKV_data_out_20_15,
           QKV_data_out_21_0, QKV_data_out_21_1, QKV_data_out_21_2, QKV_data_out_21_3, QKV_data_out_21_4, QKV_data_out_21_5, QKV_data_out_21_6, QKV_data_out_21_7, QKV_data_out_21_8, QKV_data_out_21_9, QKV_data_out_21_10, QKV_data_out_21_11, QKV_data_out_21_12, QKV_data_out_21_13, QKV_data_out_21_14, QKV_data_out_21_15,
           QKV_data_out_22_0, QKV_data_out_22_1, QKV_data_out_22_2, QKV_data_out_22_3, QKV_data_out_22_4, QKV_data_out_22_5, QKV_data_out_22_6, QKV_data_out_22_7, QKV_data_out_22_8, QKV_data_out_22_9, QKV_data_out_22_10, QKV_data_out_22_11, QKV_data_out_22_12, QKV_data_out_22_13, QKV_data_out_22_14, QKV_data_out_22_15,
           QKV_data_out_23_0, QKV_data_out_23_1, QKV_data_out_23_2, QKV_data_out_23_3, QKV_data_out_23_4, QKV_data_out_23_5, QKV_data_out_23_6, QKV_data_out_23_7, QKV_data_out_23_8, QKV_data_out_23_9, QKV_data_out_23_10, QKV_data_out_23_11, QKV_data_out_23_12, QKV_data_out_23_13, QKV_data_out_23_14, QKV_data_out_23_15,
           QKV_data_out_24_0, QKV_data_out_24_1, QKV_data_out_24_2, QKV_data_out_24_3, QKV_data_out_24_4, QKV_data_out_24_5, QKV_data_out_24_6, QKV_data_out_24_7, QKV_data_out_24_8, QKV_data_out_24_9, QKV_data_out_24_10, QKV_data_out_24_11, QKV_data_out_24_12, QKV_data_out_24_13, QKV_data_out_24_14, QKV_data_out_24_15,
           QKV_data_out_25_0, QKV_data_out_25_1, QKV_data_out_25_2, QKV_data_out_25_3, QKV_data_out_25_4, QKV_data_out_25_5, QKV_data_out_25_6, QKV_data_out_25_7, QKV_data_out_25_8, QKV_data_out_25_9, QKV_data_out_25_10, QKV_data_out_25_11, QKV_data_out_25_12, QKV_data_out_25_13, QKV_data_out_25_14, QKV_data_out_25_15,
           QKV_data_out_26_0, QKV_data_out_26_1, QKV_data_out_26_2, QKV_data_out_26_3, QKV_data_out_26_4, QKV_data_out_26_5, QKV_data_out_26_6, QKV_data_out_26_7, QKV_data_out_26_8, QKV_data_out_26_9, QKV_data_out_26_10, QKV_data_out_26_11, QKV_data_out_26_12, QKV_data_out_26_13, QKV_data_out_26_14, QKV_data_out_26_15,
           QKV_data_out_27_0, QKV_data_out_27_1, QKV_data_out_27_2, QKV_data_out_27_3, QKV_data_out_27_4, QKV_data_out_27_5, QKV_data_out_27_6, QKV_data_out_27_7, QKV_data_out_27_8, QKV_data_out_27_9, QKV_data_out_27_10, QKV_data_out_27_11, QKV_data_out_27_12, QKV_data_out_27_13, QKV_data_out_27_14, QKV_data_out_27_15,
           QKV_data_out_28_0, QKV_data_out_28_1, QKV_data_out_28_2, QKV_data_out_28_3, QKV_data_out_28_4, QKV_data_out_28_5, QKV_data_out_28_6, QKV_data_out_28_7, QKV_data_out_28_8, QKV_data_out_28_9, QKV_data_out_28_10, QKV_data_out_28_11, QKV_data_out_28_12, QKV_data_out_28_13, QKV_data_out_28_14, QKV_data_out_28_15,
           QKV_data_out_29_0, QKV_data_out_29_1, QKV_data_out_29_2, QKV_data_out_29_3, QKV_data_out_29_4, QKV_data_out_29_5, QKV_data_out_29_6, QKV_data_out_29_7, QKV_data_out_29_8, QKV_data_out_29_9, QKV_data_out_29_10, QKV_data_out_29_11, QKV_data_out_29_12, QKV_data_out_29_13, QKV_data_out_29_14, QKV_data_out_29_15,
           QKV_data_out_30_0, QKV_data_out_30_1, QKV_data_out_30_2, QKV_data_out_30_3, QKV_data_out_30_4, QKV_data_out_30_5, QKV_data_out_30_6, QKV_data_out_30_7, QKV_data_out_30_8, QKV_data_out_30_9, QKV_data_out_30_10, QKV_data_out_30_11, QKV_data_out_30_12, QKV_data_out_30_13, QKV_data_out_30_14, QKV_data_out_30_15,
           QKV_data_out_31_0, QKV_data_out_31_1, QKV_data_out_31_2, QKV_data_out_31_3, QKV_data_out_31_4, QKV_data_out_31_5, QKV_data_out_31_6, QKV_data_out_31_7, QKV_data_out_31_8, QKV_data_out_31_9, QKV_data_out_31_10, QKV_data_out_31_11, QKV_data_out_31_12, QKV_data_out_31_13, QKV_data_out_31_14, QKV_data_out_31_15;

wire [3:0] QKT_data_out_0_0, QKT_data_out_0_1, QKT_data_out_0_2, QKT_data_out_0_3, QKT_data_out_0_4, QKT_data_out_0_5, QKT_data_out_0_6, QKT_data_out_0_7, QKT_data_out_0_8, QKT_data_out_0_9, QKT_data_out_0_10, QKT_data_out_0_11, QKT_data_out_0_12, QKT_data_out_0_13, QKT_data_out_0_14, QKT_data_out_0_15,
           QKT_data_out_1_0, QKT_data_out_1_1, QKT_data_out_1_2, QKT_data_out_1_3, QKT_data_out_1_4, QKT_data_out_1_5, QKT_data_out_1_6, QKT_data_out_1_7, QKT_data_out_1_8, QKT_data_out_1_9, QKT_data_out_1_10, QKT_data_out_1_11, QKT_data_out_1_12, QKT_data_out_1_13, QKT_data_out_1_14, QKT_data_out_1_15,
           QKT_data_out_2_0, QKT_data_out_2_1, QKT_data_out_2_2, QKT_data_out_2_3, QKT_data_out_2_4, QKT_data_out_2_5, QKT_data_out_2_6, QKT_data_out_2_7, QKT_data_out_2_8, QKT_data_out_2_9, QKT_data_out_2_10, QKT_data_out_2_11, QKT_data_out_2_12, QKT_data_out_2_13, QKT_data_out_2_14, QKT_data_out_2_15,
           QKT_data_out_3_0, QKT_data_out_3_1, QKT_data_out_3_2, QKT_data_out_3_3, QKT_data_out_3_4, QKT_data_out_3_5, QKT_data_out_3_6, QKT_data_out_3_7, QKT_data_out_3_8, QKT_data_out_3_9, QKT_data_out_3_10, QKT_data_out_3_11, QKT_data_out_3_12, QKT_data_out_3_13, QKT_data_out_3_14, QKT_data_out_3_15;

wire       QKV_is_write_out_0, QKV_is_write_out_1, QKV_is_write_out_2, QKV_is_write_out_3, QKV_is_write_out_4, QKV_is_write_out_5, QKV_is_write_out_6, QKV_is_write_out_7, QKV_is_write_out_8, QKV_is_write_out_9, QKV_is_write_out_10, QKV_is_write_out_11, QKV_is_write_out_12, QKV_is_write_out_13, QKV_is_write_out_14, QKV_is_write_out_15, 
           QKV_is_write_out_16, QKV_is_write_out_17, QKV_is_write_out_18, QKV_is_write_out_19, QKV_is_write_out_20, QKV_is_write_out_21, QKV_is_write_out_22, QKV_is_write_out_23, QKV_is_write_out_24, QKV_is_write_out_25, QKV_is_write_out_26, QKV_is_write_out_27, QKV_is_write_out_28, QKV_is_write_out_29, QKV_is_write_out_30, QKV_is_write_out_31;

wire       QKT_is_write_out_0, QKT_is_write_out_1, QKT_is_write_out_2, QKT_is_write_out_3;

wire       QKV_selcet_out_0, QKV_selcet_out_1, QKV_selcet_out_2, QKV_selcet_out_3, QKV_selcet_out_4, QKV_selcet_out_5, QKV_selcet_out_6, QKV_selcet_out_7, QKV_selcet_out_8, QKV_selcet_out_9, QKV_selcet_out_10, QKV_selcet_out_11, QKV_selcet_out_12, QKV_selcet_out_13, QKV_selcet_out_14, QKV_selcet_out_15, 
           QKV_selcet_out_16, QKV_selcet_out_17, QKV_selcet_out_18, QKV_selcet_out_19, QKV_selcet_out_20, QKV_selcet_out_21, QKV_selcet_out_22, QKV_selcet_out_23, QKV_selcet_out_24, QKV_selcet_out_25, QKV_selcet_out_26, QKV_selcet_out_27, QKV_selcet_out_28, QKV_selcet_out_29, QKV_selcet_out_30, QKV_selcet_out_31;

wire       QKT_select_out_0, QKT_select_out_1, QKT_select_out_2, QKT_select_out_3;

snax_interfaces i_snax_interfaces(
    .clk(clk_i),
    .rst(rst),

    .snax_acc_req_valid(csr_req_valid_i),
    .snax_acc_req_data_addr(csr_req_addr_i),
    .snax_acc_req_data_wen(csr_req_write_i),
    .snax_acc_req_data_data(csr_req_data_i),
    .snax_acc_req_ready(csr_req_ready_o),

    .acc_snax_rsp_valid(csr_rsp_valid_o),
    .acc_snax_rsp_data_data(csr_rsp_data_o),
    .acc_snax_rsp_ready(csr_rsp_ready_i),

    .stream_acc_port_0_valid(stream2acc_0_valid_i),
    .stream_acc_port_0_data(stream2acc_0_data_i),
    .stream_acc_port_0_ready(stream2acc_0_ready_o),

    .stream_acc_port_1_valid(stream2acc_1_valid_i),
    .stream_acc_port_1_data(stream2acc_1_data_i),
    .stream_acc_port_1_ready(stream2acc_1_ready_o),

    .stream_acc_port_2_valid(stream2acc_2_valid_i),
    .stream_acc_port_2_data(stream2acc_2_data_i),
    .stream_acc_port_2_ready(stream2acc_2_ready_o),

    .stream_acc_port_3_valid(stream2acc_3_valid_i),
    .stream_acc_port_3_data(stream2acc_3_data_i),
    .stream_acc_port_3_ready(stream2acc_3_ready_o),

    .acc_stream_port_valid(acc2stream_0_valid_o),
    .acc_stream_port_data(acc2stream_0_data_o),
    .acc_stream_port_ready(acc2stream_0_ready_i),

    .QKV_addr_out_0(QKV_addr_out_0), 
    .QKV_addr_out_1(QKV_addr_out_1), 
    .QKV_addr_out_2(QKV_addr_out_2), 
    .QKV_addr_out_3(QKV_addr_out_3), 
    .QKV_addr_out_4(QKV_addr_out_4), 
    .QKV_addr_out_5(QKV_addr_out_5), 
    .QKV_addr_out_6(QKV_addr_out_6), 
    .QKV_addr_out_7(QKV_addr_out_7), 
    .QKV_addr_out_8(QKV_addr_out_8), 
    .QKV_addr_out_9(QKV_addr_out_9), 

    .QKV_addr_out_10(QKV_addr_out_10),
    .QKV_addr_out_11(QKV_addr_out_11),
    .QKV_addr_out_12(QKV_addr_out_12),
    .QKV_addr_out_13(QKV_addr_out_13),
    .QKV_addr_out_14(QKV_addr_out_14),
    .QKV_addr_out_15(QKV_addr_out_15),
    .QKV_addr_out_16(QKV_addr_out_16),
    .QKV_addr_out_17(QKV_addr_out_17),
    .QKV_addr_out_18(QKV_addr_out_18),
    .QKV_addr_out_19(QKV_addr_out_19),

    .QKV_addr_out_20(QKV_addr_out_20),
    .QKV_addr_out_21(QKV_addr_out_21),
    .QKV_addr_out_22(QKV_addr_out_22),
    .QKV_addr_out_23(QKV_addr_out_23),
    .QKV_addr_out_24(QKV_addr_out_24),
    .QKV_addr_out_25(QKV_addr_out_25),
    .QKV_addr_out_26(QKV_addr_out_26),
    .QKV_addr_out_27(QKV_addr_out_27),
    .QKV_addr_out_28(QKV_addr_out_28),
    .QKV_addr_out_29(QKV_addr_out_29),

    .QKV_addr_out_30(QKV_addr_out_30),
    .QKV_addr_out_31(QKV_addr_out_31),
    
    .QKV_calc_result_0_0(QKV_calc_result_0_0), .QKV_calc_result_0_1(QKV_calc_result_0_1), .QKV_calc_result_0_2(QKV_calc_result_0_2), .QKV_calc_result_0_3(QKV_calc_result_0_3), .QKV_calc_result_0_4(QKV_calc_result_0_4), .QKV_calc_result_0_5(QKV_calc_result_0_5), .QKV_calc_result_0_6(QKV_calc_result_0_6), .QKV_calc_result_0_7(QKV_calc_result_0_7), .QKV_calc_result_0_8(QKV_calc_result_0_8), .QKV_calc_result_0_9(QKV_calc_result_0_9), .QKV_calc_result_0_10(QKV_calc_result_0_10), .QKV_calc_result_0_11(QKV_calc_result_0_11), .QKV_calc_result_0_12(QKV_calc_result_0_12), .QKV_calc_result_0_13(QKV_calc_result_0_13), .QKV_calc_result_0_14(QKV_calc_result_0_14), .QKV_calc_result_0_15(QKV_calc_result_0_15),
    .QKV_calc_result_1_0(QKV_calc_result_1_0), .QKV_calc_result_1_1(QKV_calc_result_1_1), .QKV_calc_result_1_2(QKV_calc_result_1_2), .QKV_calc_result_1_3(QKV_calc_result_1_3), .QKV_calc_result_1_4(QKV_calc_result_1_4), .QKV_calc_result_1_5(QKV_calc_result_1_5), .QKV_calc_result_1_6(QKV_calc_result_1_6), .QKV_calc_result_1_7(QKV_calc_result_1_7), .QKV_calc_result_1_8(QKV_calc_result_1_8), .QKV_calc_result_1_9(QKV_calc_result_1_9), .QKV_calc_result_1_10(QKV_calc_result_1_10), .QKV_calc_result_1_11(QKV_calc_result_1_11), .QKV_calc_result_1_12(QKV_calc_result_1_12), .QKV_calc_result_1_13(QKV_calc_result_1_13), .QKV_calc_result_1_14(QKV_calc_result_1_14), .QKV_calc_result_1_15(QKV_calc_result_1_15),
    .QKV_calc_result_2_0(QKV_calc_result_2_0), .QKV_calc_result_2_1(QKV_calc_result_2_1), .QKV_calc_result_2_2(QKV_calc_result_2_2), .QKV_calc_result_2_3(QKV_calc_result_2_3), .QKV_calc_result_2_4(QKV_calc_result_2_4), .QKV_calc_result_2_5(QKV_calc_result_2_5), .QKV_calc_result_2_6(QKV_calc_result_2_6), .QKV_calc_result_2_7(QKV_calc_result_2_7), .QKV_calc_result_2_8(QKV_calc_result_2_8), .QKV_calc_result_2_9(QKV_calc_result_2_9), .QKV_calc_result_2_10(QKV_calc_result_2_10), .QKV_calc_result_2_11(QKV_calc_result_2_11), .QKV_calc_result_2_12(QKV_calc_result_2_12), .QKV_calc_result_2_13(QKV_calc_result_2_13), .QKV_calc_result_2_14(QKV_calc_result_2_14), .QKV_calc_result_2_15(QKV_calc_result_2_15),
    .QKV_calc_result_3_0(QKV_calc_result_3_0), .QKV_calc_result_3_1(QKV_calc_result_3_1), .QKV_calc_result_3_2(QKV_calc_result_3_2), .QKV_calc_result_3_3(QKV_calc_result_3_3), .QKV_calc_result_3_4(QKV_calc_result_3_4), .QKV_calc_result_3_5(QKV_calc_result_3_5), .QKV_calc_result_3_6(QKV_calc_result_3_6), .QKV_calc_result_3_7(QKV_calc_result_3_7), .QKV_calc_result_3_8(QKV_calc_result_3_8), .QKV_calc_result_3_9(QKV_calc_result_3_9), .QKV_calc_result_3_10(QKV_calc_result_3_10), .QKV_calc_result_3_11(QKV_calc_result_3_11), .QKV_calc_result_3_12(QKV_calc_result_3_12), .QKV_calc_result_3_13(QKV_calc_result_3_13), .QKV_calc_result_3_14(QKV_calc_result_3_14), .QKV_calc_result_3_15(QKV_calc_result_3_15),
    .QKV_calc_result_4_0(QKV_calc_result_4_0), .QKV_calc_result_4_1(QKV_calc_result_4_1), .QKV_calc_result_4_2(QKV_calc_result_4_2), .QKV_calc_result_4_3(QKV_calc_result_4_3), .QKV_calc_result_4_4(QKV_calc_result_4_4), .QKV_calc_result_4_5(QKV_calc_result_4_5), .QKV_calc_result_4_6(QKV_calc_result_4_6), .QKV_calc_result_4_7(QKV_calc_result_4_7), .QKV_calc_result_4_8(QKV_calc_result_4_8), .QKV_calc_result_4_9(QKV_calc_result_4_9), .QKV_calc_result_4_10(QKV_calc_result_4_10), .QKV_calc_result_4_11(QKV_calc_result_4_11), .QKV_calc_result_4_12(QKV_calc_result_4_12), .QKV_calc_result_4_13(QKV_calc_result_4_13), .QKV_calc_result_4_14(QKV_calc_result_4_14), .QKV_calc_result_4_15(QKV_calc_result_4_15),
    .QKV_calc_result_5_0(QKV_calc_result_5_0), .QKV_calc_result_5_1(QKV_calc_result_5_1), .QKV_calc_result_5_2(QKV_calc_result_5_2), .QKV_calc_result_5_3(QKV_calc_result_5_3), .QKV_calc_result_5_4(QKV_calc_result_5_4), .QKV_calc_result_5_5(QKV_calc_result_5_5), .QKV_calc_result_5_6(QKV_calc_result_5_6), .QKV_calc_result_5_7(QKV_calc_result_5_7), .QKV_calc_result_5_8(QKV_calc_result_5_8), .QKV_calc_result_5_9(QKV_calc_result_5_9), .QKV_calc_result_5_10(QKV_calc_result_5_10), .QKV_calc_result_5_11(QKV_calc_result_5_11), .QKV_calc_result_5_12(QKV_calc_result_5_12), .QKV_calc_result_5_13(QKV_calc_result_5_13), .QKV_calc_result_5_14(QKV_calc_result_5_14), .QKV_calc_result_5_15(QKV_calc_result_5_15),
    .QKV_calc_result_6_0(QKV_calc_result_6_0), .QKV_calc_result_6_1(QKV_calc_result_6_1), .QKV_calc_result_6_2(QKV_calc_result_6_2), .QKV_calc_result_6_3(QKV_calc_result_6_3), .QKV_calc_result_6_4(QKV_calc_result_6_4), .QKV_calc_result_6_5(QKV_calc_result_6_5), .QKV_calc_result_6_6(QKV_calc_result_6_6), .QKV_calc_result_6_7(QKV_calc_result_6_7), .QKV_calc_result_6_8(QKV_calc_result_6_8), .QKV_calc_result_6_9(QKV_calc_result_6_9), .QKV_calc_result_6_10(QKV_calc_result_6_10), .QKV_calc_result_6_11(QKV_calc_result_6_11), .QKV_calc_result_6_12(QKV_calc_result_6_12), .QKV_calc_result_6_13(QKV_calc_result_6_13), .QKV_calc_result_6_14(QKV_calc_result_6_14), .QKV_calc_result_6_15(QKV_calc_result_6_15),
    .QKV_calc_result_7_0(QKV_calc_result_7_0), .QKV_calc_result_7_1(QKV_calc_result_7_1), .QKV_calc_result_7_2(QKV_calc_result_7_2), .QKV_calc_result_7_3(QKV_calc_result_7_3), .QKV_calc_result_7_4(QKV_calc_result_7_4), .QKV_calc_result_7_5(QKV_calc_result_7_5), .QKV_calc_result_7_6(QKV_calc_result_7_6), .QKV_calc_result_7_7(QKV_calc_result_7_7), .QKV_calc_result_7_8(QKV_calc_result_7_8), .QKV_calc_result_7_9(QKV_calc_result_7_9), .QKV_calc_result_7_10(QKV_calc_result_7_10), .QKV_calc_result_7_11(QKV_calc_result_7_11), .QKV_calc_result_7_12(QKV_calc_result_7_12), .QKV_calc_result_7_13(QKV_calc_result_7_13), .QKV_calc_result_7_14(QKV_calc_result_7_14), .QKV_calc_result_7_15(QKV_calc_result_7_15),
    .QKV_calc_result_8_0(QKV_calc_result_8_0), .QKV_calc_result_8_1(QKV_calc_result_8_1), .QKV_calc_result_8_2(QKV_calc_result_8_2), .QKV_calc_result_8_3(QKV_calc_result_8_3), .QKV_calc_result_8_4(QKV_calc_result_8_4), .QKV_calc_result_8_5(QKV_calc_result_8_5), .QKV_calc_result_8_6(QKV_calc_result_8_6), .QKV_calc_result_8_7(QKV_calc_result_8_7), .QKV_calc_result_8_8(QKV_calc_result_8_8), .QKV_calc_result_8_9(QKV_calc_result_8_9), .QKV_calc_result_8_10(QKV_calc_result_8_10), .QKV_calc_result_8_11(QKV_calc_result_8_11), .QKV_calc_result_8_12(QKV_calc_result_8_12), .QKV_calc_result_8_13(QKV_calc_result_8_13), .QKV_calc_result_8_14(QKV_calc_result_8_14), .QKV_calc_result_8_15(QKV_calc_result_8_15),
    .QKV_calc_result_9_0(QKV_calc_result_9_0), .QKV_calc_result_9_1(QKV_calc_result_9_1), .QKV_calc_result_9_2(QKV_calc_result_9_2), .QKV_calc_result_9_3(QKV_calc_result_9_3), .QKV_calc_result_9_4(QKV_calc_result_9_4), .QKV_calc_result_9_5(QKV_calc_result_9_5), .QKV_calc_result_9_6(QKV_calc_result_9_6), .QKV_calc_result_9_7(QKV_calc_result_9_7), .QKV_calc_result_9_8(QKV_calc_result_9_8), .QKV_calc_result_9_9(QKV_calc_result_9_9), .QKV_calc_result_9_10(QKV_calc_result_9_10), .QKV_calc_result_9_11(QKV_calc_result_9_11), .QKV_calc_result_9_12(QKV_calc_result_9_12), .QKV_calc_result_9_13(QKV_calc_result_9_13), .QKV_calc_result_9_14(QKV_calc_result_9_14), .QKV_calc_result_9_15(QKV_calc_result_9_15),
    .QKV_calc_result_10_0(QKV_calc_result_10_0), .QKV_calc_result_10_1(QKV_calc_result_10_1), .QKV_calc_result_10_2(QKV_calc_result_10_2), .QKV_calc_result_10_3(QKV_calc_result_10_3), .QKV_calc_result_10_4(QKV_calc_result_10_4), .QKV_calc_result_10_5(QKV_calc_result_10_5), .QKV_calc_result_10_6(QKV_calc_result_10_6), .QKV_calc_result_10_7(QKV_calc_result_10_7), .QKV_calc_result_10_8(QKV_calc_result_10_8), .QKV_calc_result_10_9(QKV_calc_result_10_9), .QKV_calc_result_10_10(QKV_calc_result_10_10), .QKV_calc_result_10_11(QKV_calc_result_10_11), .QKV_calc_result_10_12(QKV_calc_result_10_12), .QKV_calc_result_10_13(QKV_calc_result_10_13), .QKV_calc_result_10_14(QKV_calc_result_10_14), .QKV_calc_result_10_15(QKV_calc_result_10_15),
    .QKV_calc_result_11_0(QKV_calc_result_11_0), .QKV_calc_result_11_1(QKV_calc_result_11_1), .QKV_calc_result_11_2(QKV_calc_result_11_2), .QKV_calc_result_11_3(QKV_calc_result_11_3), .QKV_calc_result_11_4(QKV_calc_result_11_4), .QKV_calc_result_11_5(QKV_calc_result_11_5), .QKV_calc_result_11_6(QKV_calc_result_11_6), .QKV_calc_result_11_7(QKV_calc_result_11_7), .QKV_calc_result_11_8(QKV_calc_result_11_8), .QKV_calc_result_11_9(QKV_calc_result_11_9), .QKV_calc_result_11_10(QKV_calc_result_11_10), .QKV_calc_result_11_11(QKV_calc_result_11_11), .QKV_calc_result_11_12(QKV_calc_result_11_12), .QKV_calc_result_11_13(QKV_calc_result_11_13), .QKV_calc_result_11_14(QKV_calc_result_11_14), .QKV_calc_result_11_15(QKV_calc_result_11_15),
    .QKV_calc_result_12_0(QKV_calc_result_12_0), .QKV_calc_result_12_1(QKV_calc_result_12_1), .QKV_calc_result_12_2(QKV_calc_result_12_2), .QKV_calc_result_12_3(QKV_calc_result_12_3), .QKV_calc_result_12_4(QKV_calc_result_12_4), .QKV_calc_result_12_5(QKV_calc_result_12_5), .QKV_calc_result_12_6(QKV_calc_result_12_6), .QKV_calc_result_12_7(QKV_calc_result_12_7), .QKV_calc_result_12_8(QKV_calc_result_12_8), .QKV_calc_result_12_9(QKV_calc_result_12_9), .QKV_calc_result_12_10(QKV_calc_result_12_10), .QKV_calc_result_12_11(QKV_calc_result_12_11), .QKV_calc_result_12_12(QKV_calc_result_12_12), .QKV_calc_result_12_13(QKV_calc_result_12_13), .QKV_calc_result_12_14(QKV_calc_result_12_14), .QKV_calc_result_12_15(QKV_calc_result_12_15),
    .QKV_calc_result_13_0(QKV_calc_result_13_0), .QKV_calc_result_13_1(QKV_calc_result_13_1), .QKV_calc_result_13_2(QKV_calc_result_13_2), .QKV_calc_result_13_3(QKV_calc_result_13_3), .QKV_calc_result_13_4(QKV_calc_result_13_4), .QKV_calc_result_13_5(QKV_calc_result_13_5), .QKV_calc_result_13_6(QKV_calc_result_13_6), .QKV_calc_result_13_7(QKV_calc_result_13_7), .QKV_calc_result_13_8(QKV_calc_result_13_8), .QKV_calc_result_13_9(QKV_calc_result_13_9), .QKV_calc_result_13_10(QKV_calc_result_13_10), .QKV_calc_result_13_11(QKV_calc_result_13_11), .QKV_calc_result_13_12(QKV_calc_result_13_12), .QKV_calc_result_13_13(QKV_calc_result_13_13), .QKV_calc_result_13_14(QKV_calc_result_13_14), .QKV_calc_result_13_15(QKV_calc_result_13_15),
    .QKV_calc_result_14_0(QKV_calc_result_14_0), .QKV_calc_result_14_1(QKV_calc_result_14_1), .QKV_calc_result_14_2(QKV_calc_result_14_2), .QKV_calc_result_14_3(QKV_calc_result_14_3), .QKV_calc_result_14_4(QKV_calc_result_14_4), .QKV_calc_result_14_5(QKV_calc_result_14_5), .QKV_calc_result_14_6(QKV_calc_result_14_6), .QKV_calc_result_14_7(QKV_calc_result_14_7), .QKV_calc_result_14_8(QKV_calc_result_14_8), .QKV_calc_result_14_9(QKV_calc_result_14_9), .QKV_calc_result_14_10(QKV_calc_result_14_10), .QKV_calc_result_14_11(QKV_calc_result_14_11), .QKV_calc_result_14_12(QKV_calc_result_14_12), .QKV_calc_result_14_13(QKV_calc_result_14_13), .QKV_calc_result_14_14(QKV_calc_result_14_14), .QKV_calc_result_14_15(QKV_calc_result_14_15),
    .QKV_calc_result_15_0(QKV_calc_result_15_0), .QKV_calc_result_15_1(QKV_calc_result_15_1), .QKV_calc_result_15_2(QKV_calc_result_15_2), .QKV_calc_result_15_3(QKV_calc_result_15_3), .QKV_calc_result_15_4(QKV_calc_result_15_4), .QKV_calc_result_15_5(QKV_calc_result_15_5), .QKV_calc_result_15_6(QKV_calc_result_15_6), .QKV_calc_result_15_7(QKV_calc_result_15_7), .QKV_calc_result_15_8(QKV_calc_result_15_8), .QKV_calc_result_15_9(QKV_calc_result_15_9), .QKV_calc_result_15_10(QKV_calc_result_15_10), .QKV_calc_result_15_11(QKV_calc_result_15_11), .QKV_calc_result_15_12(QKV_calc_result_15_12), .QKV_calc_result_15_13(QKV_calc_result_15_13), .QKV_calc_result_15_14(QKV_calc_result_15_14), .QKV_calc_result_15_15(QKV_calc_result_15_15),
    .QKV_calc_result_16_0(QKV_calc_result_16_0), .QKV_calc_result_16_1(QKV_calc_result_16_1), .QKV_calc_result_16_2(QKV_calc_result_16_2), .QKV_calc_result_16_3(QKV_calc_result_16_3), .QKV_calc_result_16_4(QKV_calc_result_16_4), .QKV_calc_result_16_5(QKV_calc_result_16_5), .QKV_calc_result_16_6(QKV_calc_result_16_6), .QKV_calc_result_16_7(QKV_calc_result_16_7), .QKV_calc_result_16_8(QKV_calc_result_16_8), .QKV_calc_result_16_9(QKV_calc_result_16_9), .QKV_calc_result_16_10(QKV_calc_result_16_10), .QKV_calc_result_16_11(QKV_calc_result_16_11), .QKV_calc_result_16_12(QKV_calc_result_16_12), .QKV_calc_result_16_13(QKV_calc_result_16_13), .QKV_calc_result_16_14(QKV_calc_result_16_14), .QKV_calc_result_16_15(QKV_calc_result_16_15),
    .QKV_calc_result_17_0(QKV_calc_result_17_0), .QKV_calc_result_17_1(QKV_calc_result_17_1), .QKV_calc_result_17_2(QKV_calc_result_17_2), .QKV_calc_result_17_3(QKV_calc_result_17_3), .QKV_calc_result_17_4(QKV_calc_result_17_4), .QKV_calc_result_17_5(QKV_calc_result_17_5), .QKV_calc_result_17_6(QKV_calc_result_17_6), .QKV_calc_result_17_7(QKV_calc_result_17_7), .QKV_calc_result_17_8(QKV_calc_result_17_8), .QKV_calc_result_17_9(QKV_calc_result_17_9), .QKV_calc_result_17_10(QKV_calc_result_17_10), .QKV_calc_result_17_11(QKV_calc_result_17_11), .QKV_calc_result_17_12(QKV_calc_result_17_12), .QKV_calc_result_17_13(QKV_calc_result_17_13), .QKV_calc_result_17_14(QKV_calc_result_17_14), .QKV_calc_result_17_15(QKV_calc_result_17_15),
    .QKV_calc_result_18_0(QKV_calc_result_18_0), .QKV_calc_result_18_1(QKV_calc_result_18_1), .QKV_calc_result_18_2(QKV_calc_result_18_2), .QKV_calc_result_18_3(QKV_calc_result_18_3), .QKV_calc_result_18_4(QKV_calc_result_18_4), .QKV_calc_result_18_5(QKV_calc_result_18_5), .QKV_calc_result_18_6(QKV_calc_result_18_6), .QKV_calc_result_18_7(QKV_calc_result_18_7), .QKV_calc_result_18_8(QKV_calc_result_18_8), .QKV_calc_result_18_9(QKV_calc_result_18_9), .QKV_calc_result_18_10(QKV_calc_result_18_10), .QKV_calc_result_18_11(QKV_calc_result_18_11), .QKV_calc_result_18_12(QKV_calc_result_18_12), .QKV_calc_result_18_13(QKV_calc_result_18_13), .QKV_calc_result_18_14(QKV_calc_result_18_14), .QKV_calc_result_18_15(QKV_calc_result_18_15),
    .QKV_calc_result_19_0(QKV_calc_result_19_0), .QKV_calc_result_19_1(QKV_calc_result_19_1), .QKV_calc_result_19_2(QKV_calc_result_19_2), .QKV_calc_result_19_3(QKV_calc_result_19_3), .QKV_calc_result_19_4(QKV_calc_result_19_4), .QKV_calc_result_19_5(QKV_calc_result_19_5), .QKV_calc_result_19_6(QKV_calc_result_19_6), .QKV_calc_result_19_7(QKV_calc_result_19_7), .QKV_calc_result_19_8(QKV_calc_result_19_8), .QKV_calc_result_19_9(QKV_calc_result_19_9), .QKV_calc_result_19_10(QKV_calc_result_19_10), .QKV_calc_result_19_11(QKV_calc_result_19_11), .QKV_calc_result_19_12(QKV_calc_result_19_12), .QKV_calc_result_19_13(QKV_calc_result_19_13), .QKV_calc_result_19_14(QKV_calc_result_19_14), .QKV_calc_result_19_15(QKV_calc_result_19_15),
    .QKV_calc_result_20_0(QKV_calc_result_20_0), .QKV_calc_result_20_1(QKV_calc_result_20_1), .QKV_calc_result_20_2(QKV_calc_result_20_2), .QKV_calc_result_20_3(QKV_calc_result_20_3), .QKV_calc_result_20_4(QKV_calc_result_20_4), .QKV_calc_result_20_5(QKV_calc_result_20_5), .QKV_calc_result_20_6(QKV_calc_result_20_6), .QKV_calc_result_20_7(QKV_calc_result_20_7), .QKV_calc_result_20_8(QKV_calc_result_20_8), .QKV_calc_result_20_9(QKV_calc_result_20_9), .QKV_calc_result_20_10(QKV_calc_result_20_10), .QKV_calc_result_20_11(QKV_calc_result_20_11), .QKV_calc_result_20_12(QKV_calc_result_20_12), .QKV_calc_result_20_13(QKV_calc_result_20_13), .QKV_calc_result_20_14(QKV_calc_result_20_14), .QKV_calc_result_20_15(QKV_calc_result_20_15),
    .QKV_calc_result_21_0(QKV_calc_result_21_0), .QKV_calc_result_21_1(QKV_calc_result_21_1), .QKV_calc_result_21_2(QKV_calc_result_21_2), .QKV_calc_result_21_3(QKV_calc_result_21_3), .QKV_calc_result_21_4(QKV_calc_result_21_4), .QKV_calc_result_21_5(QKV_calc_result_21_5), .QKV_calc_result_21_6(QKV_calc_result_21_6), .QKV_calc_result_21_7(QKV_calc_result_21_7), .QKV_calc_result_21_8(QKV_calc_result_21_8), .QKV_calc_result_21_9(QKV_calc_result_21_9), .QKV_calc_result_21_10(QKV_calc_result_21_10), .QKV_calc_result_21_11(QKV_calc_result_21_11), .QKV_calc_result_21_12(QKV_calc_result_21_12), .QKV_calc_result_21_13(QKV_calc_result_21_13), .QKV_calc_result_21_14(QKV_calc_result_21_14), .QKV_calc_result_21_15(QKV_calc_result_21_15),
    .QKV_calc_result_22_0(QKV_calc_result_22_0), .QKV_calc_result_22_1(QKV_calc_result_22_1), .QKV_calc_result_22_2(QKV_calc_result_22_2), .QKV_calc_result_22_3(QKV_calc_result_22_3), .QKV_calc_result_22_4(QKV_calc_result_22_4), .QKV_calc_result_22_5(QKV_calc_result_22_5), .QKV_calc_result_22_6(QKV_calc_result_22_6), .QKV_calc_result_22_7(QKV_calc_result_22_7), .QKV_calc_result_22_8(QKV_calc_result_22_8), .QKV_calc_result_22_9(QKV_calc_result_22_9), .QKV_calc_result_22_10(QKV_calc_result_22_10), .QKV_calc_result_22_11(QKV_calc_result_22_11), .QKV_calc_result_22_12(QKV_calc_result_22_12), .QKV_calc_result_22_13(QKV_calc_result_22_13), .QKV_calc_result_22_14(QKV_calc_result_22_14), .QKV_calc_result_22_15(QKV_calc_result_22_15),
    .QKV_calc_result_23_0(QKV_calc_result_23_0), .QKV_calc_result_23_1(QKV_calc_result_23_1), .QKV_calc_result_23_2(QKV_calc_result_23_2), .QKV_calc_result_23_3(QKV_calc_result_23_3), .QKV_calc_result_23_4(QKV_calc_result_23_4), .QKV_calc_result_23_5(QKV_calc_result_23_5), .QKV_calc_result_23_6(QKV_calc_result_23_6), .QKV_calc_result_23_7(QKV_calc_result_23_7), .QKV_calc_result_23_8(QKV_calc_result_23_8), .QKV_calc_result_23_9(QKV_calc_result_23_9), .QKV_calc_result_23_10(QKV_calc_result_23_10), .QKV_calc_result_23_11(QKV_calc_result_23_11), .QKV_calc_result_23_12(QKV_calc_result_23_12), .QKV_calc_result_23_13(QKV_calc_result_23_13), .QKV_calc_result_23_14(QKV_calc_result_23_14), .QKV_calc_result_23_15(QKV_calc_result_23_15),
    .QKV_calc_result_24_0(QKV_calc_result_24_0), .QKV_calc_result_24_1(QKV_calc_result_24_1), .QKV_calc_result_24_2(QKV_calc_result_24_2), .QKV_calc_result_24_3(QKV_calc_result_24_3), .QKV_calc_result_24_4(QKV_calc_result_24_4), .QKV_calc_result_24_5(QKV_calc_result_24_5), .QKV_calc_result_24_6(QKV_calc_result_24_6), .QKV_calc_result_24_7(QKV_calc_result_24_7), .QKV_calc_result_24_8(QKV_calc_result_24_8), .QKV_calc_result_24_9(QKV_calc_result_24_9), .QKV_calc_result_24_10(QKV_calc_result_24_10), .QKV_calc_result_24_11(QKV_calc_result_24_11), .QKV_calc_result_24_12(QKV_calc_result_24_12), .QKV_calc_result_24_13(QKV_calc_result_24_13), .QKV_calc_result_24_14(QKV_calc_result_24_14), .QKV_calc_result_24_15(QKV_calc_result_24_15),
    .QKV_calc_result_25_0(QKV_calc_result_25_0), .QKV_calc_result_25_1(QKV_calc_result_25_1), .QKV_calc_result_25_2(QKV_calc_result_25_2), .QKV_calc_result_25_3(QKV_calc_result_25_3), .QKV_calc_result_25_4(QKV_calc_result_25_4), .QKV_calc_result_25_5(QKV_calc_result_25_5), .QKV_calc_result_25_6(QKV_calc_result_25_6), .QKV_calc_result_25_7(QKV_calc_result_25_7), .QKV_calc_result_25_8(QKV_calc_result_25_8), .QKV_calc_result_25_9(QKV_calc_result_25_9), .QKV_calc_result_25_10(QKV_calc_result_25_10), .QKV_calc_result_25_11(QKV_calc_result_25_11), .QKV_calc_result_25_12(QKV_calc_result_25_12), .QKV_calc_result_25_13(QKV_calc_result_25_13), .QKV_calc_result_25_14(QKV_calc_result_25_14), .QKV_calc_result_25_15(QKV_calc_result_25_15),
    .QKV_calc_result_26_0(QKV_calc_result_26_0), .QKV_calc_result_26_1(QKV_calc_result_26_1), .QKV_calc_result_26_2(QKV_calc_result_26_2), .QKV_calc_result_26_3(QKV_calc_result_26_3), .QKV_calc_result_26_4(QKV_calc_result_26_4), .QKV_calc_result_26_5(QKV_calc_result_26_5), .QKV_calc_result_26_6(QKV_calc_result_26_6), .QKV_calc_result_26_7(QKV_calc_result_26_7), .QKV_calc_result_26_8(QKV_calc_result_26_8), .QKV_calc_result_26_9(QKV_calc_result_26_9), .QKV_calc_result_26_10(QKV_calc_result_26_10), .QKV_calc_result_26_11(QKV_calc_result_26_11), .QKV_calc_result_26_12(QKV_calc_result_26_12), .QKV_calc_result_26_13(QKV_calc_result_26_13), .QKV_calc_result_26_14(QKV_calc_result_26_14), .QKV_calc_result_26_15(QKV_calc_result_26_15),
    .QKV_calc_result_27_0(QKV_calc_result_27_0), .QKV_calc_result_27_1(QKV_calc_result_27_1), .QKV_calc_result_27_2(QKV_calc_result_27_2), .QKV_calc_result_27_3(QKV_calc_result_27_3), .QKV_calc_result_27_4(QKV_calc_result_27_4), .QKV_calc_result_27_5(QKV_calc_result_27_5), .QKV_calc_result_27_6(QKV_calc_result_27_6), .QKV_calc_result_27_7(QKV_calc_result_27_7), .QKV_calc_result_27_8(QKV_calc_result_27_8), .QKV_calc_result_27_9(QKV_calc_result_27_9), .QKV_calc_result_27_10(QKV_calc_result_27_10), .QKV_calc_result_27_11(QKV_calc_result_27_11), .QKV_calc_result_27_12(QKV_calc_result_27_12), .QKV_calc_result_27_13(QKV_calc_result_27_13), .QKV_calc_result_27_14(QKV_calc_result_27_14), .QKV_calc_result_27_15(QKV_calc_result_27_15),
    .QKV_calc_result_28_0(QKV_calc_result_28_0), .QKV_calc_result_28_1(QKV_calc_result_28_1), .QKV_calc_result_28_2(QKV_calc_result_28_2), .QKV_calc_result_28_3(QKV_calc_result_28_3), .QKV_calc_result_28_4(QKV_calc_result_28_4), .QKV_calc_result_28_5(QKV_calc_result_28_5), .QKV_calc_result_28_6(QKV_calc_result_28_6), .QKV_calc_result_28_7(QKV_calc_result_28_7), .QKV_calc_result_28_8(QKV_calc_result_28_8), .QKV_calc_result_28_9(QKV_calc_result_28_9), .QKV_calc_result_28_10(QKV_calc_result_28_10), .QKV_calc_result_28_11(QKV_calc_result_28_11), .QKV_calc_result_28_12(QKV_calc_result_28_12), .QKV_calc_result_28_13(QKV_calc_result_28_13), .QKV_calc_result_28_14(QKV_calc_result_28_14), .QKV_calc_result_28_15(QKV_calc_result_28_15),
    .QKV_calc_result_29_0(QKV_calc_result_29_0), .QKV_calc_result_29_1(QKV_calc_result_29_1), .QKV_calc_result_29_2(QKV_calc_result_29_2), .QKV_calc_result_29_3(QKV_calc_result_29_3), .QKV_calc_result_29_4(QKV_calc_result_29_4), .QKV_calc_result_29_5(QKV_calc_result_29_5), .QKV_calc_result_29_6(QKV_calc_result_29_6), .QKV_calc_result_29_7(QKV_calc_result_29_7), .QKV_calc_result_29_8(QKV_calc_result_29_8), .QKV_calc_result_29_9(QKV_calc_result_29_9), .QKV_calc_result_29_10(QKV_calc_result_29_10), .QKV_calc_result_29_11(QKV_calc_result_29_11), .QKV_calc_result_29_12(QKV_calc_result_29_12), .QKV_calc_result_29_13(QKV_calc_result_29_13), .QKV_calc_result_29_14(QKV_calc_result_29_14), .QKV_calc_result_29_15(QKV_calc_result_29_15),
    .QKV_calc_result_30_0(QKV_calc_result_30_0), .QKV_calc_result_30_1(QKV_calc_result_30_1), .QKV_calc_result_30_2(QKV_calc_result_30_2), .QKV_calc_result_30_3(QKV_calc_result_30_3), .QKV_calc_result_30_4(QKV_calc_result_30_4), .QKV_calc_result_30_5(QKV_calc_result_30_5), .QKV_calc_result_30_6(QKV_calc_result_30_6), .QKV_calc_result_30_7(QKV_calc_result_30_7), .QKV_calc_result_30_8(QKV_calc_result_30_8), .QKV_calc_result_30_9(QKV_calc_result_30_9), .QKV_calc_result_30_10(QKV_calc_result_30_10), .QKV_calc_result_30_11(QKV_calc_result_30_11), .QKV_calc_result_30_12(QKV_calc_result_30_12), .QKV_calc_result_30_13(QKV_calc_result_30_13), .QKV_calc_result_30_14(QKV_calc_result_30_14), .QKV_calc_result_30_15(QKV_calc_result_30_15),
    .QKV_calc_result_31_0(QKV_calc_result_31_0), .QKV_calc_result_31_1(QKV_calc_result_31_1), .QKV_calc_result_31_2(QKV_calc_result_31_2), .QKV_calc_result_31_3(QKV_calc_result_31_3), .QKV_calc_result_31_4(QKV_calc_result_31_4), .QKV_calc_result_31_5(QKV_calc_result_31_5), .QKV_calc_result_31_6(QKV_calc_result_31_6), .QKV_calc_result_31_7(QKV_calc_result_31_7), .QKV_calc_result_31_8(QKV_calc_result_31_8), .QKV_calc_result_31_9(QKV_calc_result_31_9), .QKV_calc_result_31_10(QKV_calc_result_31_10), .QKV_calc_result_31_11(QKV_calc_result_31_11), .QKV_calc_result_31_12(QKV_calc_result_31_12), .QKV_calc_result_31_13(QKV_calc_result_31_13), .QKV_calc_result_31_14(QKV_calc_result_31_14), .QKV_calc_result_31_15(QKV_calc_result_31_15),

    .QKT_calc_result_0_0(QKT_calc_result_0_0), .QKT_calc_result_0_1(QKT_calc_result_0_1), .QKT_calc_result_0_2(QKT_calc_result_0_2), .QKT_calc_result_0_3(QKT_calc_result_0_3), .QKT_calc_result_0_4(QKT_calc_result_0_4), .QKT_calc_result_0_5(QKT_calc_result_0_5), .QKT_calc_result_0_6(QKT_calc_result_0_6), .QKT_calc_result_0_7(QKT_calc_result_0_7), .QKT_calc_result_0_8(QKT_calc_result_0_8), .QKT_calc_result_0_9(QKT_calc_result_0_9), .QKT_calc_result_0_10(QKT_calc_result_0_10), .QKT_calc_result_0_11(QKT_calc_result_0_11), .QKT_calc_result_0_12(QKT_calc_result_0_12), .QKT_calc_result_0_13(QKT_calc_result_0_13), .QKT_calc_result_0_14(QKT_calc_result_0_14), .QKT_calc_result_0_15(QKT_calc_result_0_15),
    .QKT_calc_result_1_0(QKT_calc_result_1_0), .QKT_calc_result_1_1(QKT_calc_result_1_1), .QKT_calc_result_1_2(QKT_calc_result_1_2), .QKT_calc_result_1_3(QKT_calc_result_1_3), .QKT_calc_result_1_4(QKT_calc_result_1_4), .QKT_calc_result_1_5(QKT_calc_result_1_5), .QKT_calc_result_1_6(QKT_calc_result_1_6), .QKT_calc_result_1_7(QKT_calc_result_1_7), .QKT_calc_result_1_8(QKT_calc_result_1_8), .QKT_calc_result_1_9(QKT_calc_result_1_9), .QKT_calc_result_1_10(QKT_calc_result_1_10), .QKT_calc_result_1_11(QKT_calc_result_1_11), .QKT_calc_result_1_12(QKT_calc_result_1_12), .QKT_calc_result_1_13(QKT_calc_result_1_13), .QKT_calc_result_1_14(QKT_calc_result_1_14), .QKT_calc_result_1_15(QKT_calc_result_1_15),
    .QKT_calc_result_2_0(QKT_calc_result_2_0), .QKT_calc_result_2_1(QKT_calc_result_2_1), .QKT_calc_result_2_2(QKT_calc_result_2_2), .QKT_calc_result_2_3(QKT_calc_result_2_3), .QKT_calc_result_2_4(QKT_calc_result_2_4), .QKT_calc_result_2_5(QKT_calc_result_2_5), .QKT_calc_result_2_6(QKT_calc_result_2_6), .QKT_calc_result_2_7(QKT_calc_result_2_7), .QKT_calc_result_2_8(QKT_calc_result_2_8), .QKT_calc_result_2_9(QKT_calc_result_2_9), .QKT_calc_result_2_10(QKT_calc_result_2_10), .QKT_calc_result_2_11(QKT_calc_result_2_11), .QKT_calc_result_2_12(QKT_calc_result_2_12), .QKT_calc_result_2_13(QKT_calc_result_2_13), .QKT_calc_result_2_14(QKT_calc_result_2_14), .QKT_calc_result_2_15(QKT_calc_result_2_15),
    .QKT_calc_result_3_0(QKT_calc_result_3_0), .QKT_calc_result_3_1(QKT_calc_result_3_1), .QKT_calc_result_3_2(QKT_calc_result_3_2), .QKT_calc_result_3_3(QKT_calc_result_3_3), .QKT_calc_result_3_4(QKT_calc_result_3_4), .QKT_calc_result_3_5(QKT_calc_result_3_5), .QKT_calc_result_3_6(QKT_calc_result_3_6), .QKT_calc_result_3_7(QKT_calc_result_3_7), .QKT_calc_result_3_8(QKT_calc_result_3_8), .QKT_calc_result_3_9(QKT_calc_result_3_9), .QKT_calc_result_3_10(QKT_calc_result_3_10), .QKT_calc_result_3_11(QKT_calc_result_3_11), .QKT_calc_result_3_12(QKT_calc_result_3_12), .QKT_calc_result_3_13(QKT_calc_result_3_13), .QKT_calc_result_3_14(QKT_calc_result_3_14), .QKT_calc_result_3_15(QKT_calc_result_3_15),

    .QKV_weight_out_0_0(QKV_weight_out_0_0), .QKV_weight_out_0_1(QKV_weight_out_0_1), .QKV_weight_out_0_2(QKV_weight_out_0_2), .QKV_weight_out_0_3(QKV_weight_out_0_3), .QKV_weight_out_0_4(QKV_weight_out_0_4), .QKV_weight_out_0_5(QKV_weight_out_0_5), .QKV_weight_out_0_6(QKV_weight_out_0_6), .QKV_weight_out_0_7(QKV_weight_out_0_7), .QKV_weight_out_0_8(QKV_weight_out_0_8), .QKV_weight_out_0_9(QKV_weight_out_0_9), .QKV_weight_out_0_10(QKV_weight_out_0_10), .QKV_weight_out_0_11(QKV_weight_out_0_11), .QKV_weight_out_0_12(QKV_weight_out_0_12), .QKV_weight_out_0_13(QKV_weight_out_0_13), .QKV_weight_out_0_14(QKV_weight_out_0_14), .QKV_weight_out_0_15(QKV_weight_out_0_15),
    .QKV_weight_out_1_0(QKV_weight_out_1_0), .QKV_weight_out_1_1(QKV_weight_out_1_1), .QKV_weight_out_1_2(QKV_weight_out_1_2), .QKV_weight_out_1_3(QKV_weight_out_1_3), .QKV_weight_out_1_4(QKV_weight_out_1_4), .QKV_weight_out_1_5(QKV_weight_out_1_5), .QKV_weight_out_1_6(QKV_weight_out_1_6), .QKV_weight_out_1_7(QKV_weight_out_1_7), .QKV_weight_out_1_8(QKV_weight_out_1_8), .QKV_weight_out_1_9(QKV_weight_out_1_9), .QKV_weight_out_1_10(QKV_weight_out_1_10), .QKV_weight_out_1_11(QKV_weight_out_1_11), .QKV_weight_out_1_12(QKV_weight_out_1_12), .QKV_weight_out_1_13(QKV_weight_out_1_13), .QKV_weight_out_1_14(QKV_weight_out_1_14), .QKV_weight_out_1_15(QKV_weight_out_1_15),
    .QKV_weight_out_2_0(QKV_weight_out_2_0), .QKV_weight_out_2_1(QKV_weight_out_2_1), .QKV_weight_out_2_2(QKV_weight_out_2_2), .QKV_weight_out_2_3(QKV_weight_out_2_3), .QKV_weight_out_2_4(QKV_weight_out_2_4), .QKV_weight_out_2_5(QKV_weight_out_2_5), .QKV_weight_out_2_6(QKV_weight_out_2_6), .QKV_weight_out_2_7(QKV_weight_out_2_7), .QKV_weight_out_2_8(QKV_weight_out_2_8), .QKV_weight_out_2_9(QKV_weight_out_2_9), .QKV_weight_out_2_10(QKV_weight_out_2_10), .QKV_weight_out_2_11(QKV_weight_out_2_11), .QKV_weight_out_2_12(QKV_weight_out_2_12), .QKV_weight_out_2_13(QKV_weight_out_2_13), .QKV_weight_out_2_14(QKV_weight_out_2_14), .QKV_weight_out_2_15(QKV_weight_out_2_15),
    .QKV_weight_out_3_0(QKV_weight_out_3_0), .QKV_weight_out_3_1(QKV_weight_out_3_1), .QKV_weight_out_3_2(QKV_weight_out_3_2), .QKV_weight_out_3_3(QKV_weight_out_3_3), .QKV_weight_out_3_4(QKV_weight_out_3_4), .QKV_weight_out_3_5(QKV_weight_out_3_5), .QKV_weight_out_3_6(QKV_weight_out_3_6), .QKV_weight_out_3_7(QKV_weight_out_3_7), .QKV_weight_out_3_8(QKV_weight_out_3_8), .QKV_weight_out_3_9(QKV_weight_out_3_9), .QKV_weight_out_3_10(QKV_weight_out_3_10), .QKV_weight_out_3_11(QKV_weight_out_3_11), .QKV_weight_out_3_12(QKV_weight_out_3_12), .QKV_weight_out_3_13(QKV_weight_out_3_13), .QKV_weight_out_3_14(QKV_weight_out_3_14), .QKV_weight_out_3_15(QKV_weight_out_3_15),
    .QKV_weight_out_4_0(QKV_weight_out_4_0), .QKV_weight_out_4_1(QKV_weight_out_4_1), .QKV_weight_out_4_2(QKV_weight_out_4_2), .QKV_weight_out_4_3(QKV_weight_out_4_3), .QKV_weight_out_4_4(QKV_weight_out_4_4), .QKV_weight_out_4_5(QKV_weight_out_4_5), .QKV_weight_out_4_6(QKV_weight_out_4_6), .QKV_weight_out_4_7(QKV_weight_out_4_7), .QKV_weight_out_4_8(QKV_weight_out_4_8), .QKV_weight_out_4_9(QKV_weight_out_4_9), .QKV_weight_out_4_10(QKV_weight_out_4_10), .QKV_weight_out_4_11(QKV_weight_out_4_11), .QKV_weight_out_4_12(QKV_weight_out_4_12), .QKV_weight_out_4_13(QKV_weight_out_4_13), .QKV_weight_out_4_14(QKV_weight_out_4_14), .QKV_weight_out_4_15(QKV_weight_out_4_15),
    .QKV_weight_out_5_0(QKV_weight_out_5_0), .QKV_weight_out_5_1(QKV_weight_out_5_1), .QKV_weight_out_5_2(QKV_weight_out_5_2), .QKV_weight_out_5_3(QKV_weight_out_5_3), .QKV_weight_out_5_4(QKV_weight_out_5_4), .QKV_weight_out_5_5(QKV_weight_out_5_5), .QKV_weight_out_5_6(QKV_weight_out_5_6), .QKV_weight_out_5_7(QKV_weight_out_5_7), .QKV_weight_out_5_8(QKV_weight_out_5_8), .QKV_weight_out_5_9(QKV_weight_out_5_9), .QKV_weight_out_5_10(QKV_weight_out_5_10), .QKV_weight_out_5_11(QKV_weight_out_5_11), .QKV_weight_out_5_12(QKV_weight_out_5_12), .QKV_weight_out_5_13(QKV_weight_out_5_13), .QKV_weight_out_5_14(QKV_weight_out_5_14), .QKV_weight_out_5_15(QKV_weight_out_5_15),
    .QKV_weight_out_6_0(QKV_weight_out_6_0), .QKV_weight_out_6_1(QKV_weight_out_6_1), .QKV_weight_out_6_2(QKV_weight_out_6_2), .QKV_weight_out_6_3(QKV_weight_out_6_3), .QKV_weight_out_6_4(QKV_weight_out_6_4), .QKV_weight_out_6_5(QKV_weight_out_6_5), .QKV_weight_out_6_6(QKV_weight_out_6_6), .QKV_weight_out_6_7(QKV_weight_out_6_7), .QKV_weight_out_6_8(QKV_weight_out_6_8), .QKV_weight_out_6_9(QKV_weight_out_6_9), .QKV_weight_out_6_10(QKV_weight_out_6_10), .QKV_weight_out_6_11(QKV_weight_out_6_11), .QKV_weight_out_6_12(QKV_weight_out_6_12), .QKV_weight_out_6_13(QKV_weight_out_6_13), .QKV_weight_out_6_14(QKV_weight_out_6_14), .QKV_weight_out_6_15(QKV_weight_out_6_15),
    .QKV_weight_out_7_0(QKV_weight_out_7_0), .QKV_weight_out_7_1(QKV_weight_out_7_1), .QKV_weight_out_7_2(QKV_weight_out_7_2), .QKV_weight_out_7_3(QKV_weight_out_7_3), .QKV_weight_out_7_4(QKV_weight_out_7_4), .QKV_weight_out_7_5(QKV_weight_out_7_5), .QKV_weight_out_7_6(QKV_weight_out_7_6), .QKV_weight_out_7_7(QKV_weight_out_7_7), .QKV_weight_out_7_8(QKV_weight_out_7_8), .QKV_weight_out_7_9(QKV_weight_out_7_9), .QKV_weight_out_7_10(QKV_weight_out_7_10), .QKV_weight_out_7_11(QKV_weight_out_7_11), .QKV_weight_out_7_12(QKV_weight_out_7_12), .QKV_weight_out_7_13(QKV_weight_out_7_13), .QKV_weight_out_7_14(QKV_weight_out_7_14), .QKV_weight_out_7_15(QKV_weight_out_7_15),
    .QKV_weight_out_8_0(QKV_weight_out_8_0), .QKV_weight_out_8_1(QKV_weight_out_8_1), .QKV_weight_out_8_2(QKV_weight_out_8_2), .QKV_weight_out_8_3(QKV_weight_out_8_3), .QKV_weight_out_8_4(QKV_weight_out_8_4), .QKV_weight_out_8_5(QKV_weight_out_8_5), .QKV_weight_out_8_6(QKV_weight_out_8_6), .QKV_weight_out_8_7(QKV_weight_out_8_7), .QKV_weight_out_8_8(QKV_weight_out_8_8), .QKV_weight_out_8_9(QKV_weight_out_8_9), .QKV_weight_out_8_10(QKV_weight_out_8_10), .QKV_weight_out_8_11(QKV_weight_out_8_11), .QKV_weight_out_8_12(QKV_weight_out_8_12), .QKV_weight_out_8_13(QKV_weight_out_8_13), .QKV_weight_out_8_14(QKV_weight_out_8_14), .QKV_weight_out_8_15(QKV_weight_out_8_15),
    .QKV_weight_out_9_0(QKV_weight_out_9_0), .QKV_weight_out_9_1(QKV_weight_out_9_1), .QKV_weight_out_9_2(QKV_weight_out_9_2), .QKV_weight_out_9_3(QKV_weight_out_9_3), .QKV_weight_out_9_4(QKV_weight_out_9_4), .QKV_weight_out_9_5(QKV_weight_out_9_5), .QKV_weight_out_9_6(QKV_weight_out_9_6), .QKV_weight_out_9_7(QKV_weight_out_9_7), .QKV_weight_out_9_8(QKV_weight_out_9_8), .QKV_weight_out_9_9(QKV_weight_out_9_9), .QKV_weight_out_9_10(QKV_weight_out_9_10), .QKV_weight_out_9_11(QKV_weight_out_9_11), .QKV_weight_out_9_12(QKV_weight_out_9_12), .QKV_weight_out_9_13(QKV_weight_out_9_13), .QKV_weight_out_9_14(QKV_weight_out_9_14), .QKV_weight_out_9_15(QKV_weight_out_9_15),
    .QKV_weight_out_10_0(QKV_weight_out_10_0), .QKV_weight_out_10_1(QKV_weight_out_10_1), .QKV_weight_out_10_2(QKV_weight_out_10_2), .QKV_weight_out_10_3(QKV_weight_out_10_3), .QKV_weight_out_10_4(QKV_weight_out_10_4), .QKV_weight_out_10_5(QKV_weight_out_10_5), .QKV_weight_out_10_6(QKV_weight_out_10_6), .QKV_weight_out_10_7(QKV_weight_out_10_7), .QKV_weight_out_10_8(QKV_weight_out_10_8), .QKV_weight_out_10_9(QKV_weight_out_10_9), .QKV_weight_out_10_10(QKV_weight_out_10_10), .QKV_weight_out_10_11(QKV_weight_out_10_11), .QKV_weight_out_10_12(QKV_weight_out_10_12), .QKV_weight_out_10_13(QKV_weight_out_10_13), .QKV_weight_out_10_14(QKV_weight_out_10_14), .QKV_weight_out_10_15(QKV_weight_out_10_15),
    .QKV_weight_out_11_0(QKV_weight_out_11_0), .QKV_weight_out_11_1(QKV_weight_out_11_1), .QKV_weight_out_11_2(QKV_weight_out_11_2), .QKV_weight_out_11_3(QKV_weight_out_11_3), .QKV_weight_out_11_4(QKV_weight_out_11_4), .QKV_weight_out_11_5(QKV_weight_out_11_5), .QKV_weight_out_11_6(QKV_weight_out_11_6), .QKV_weight_out_11_7(QKV_weight_out_11_7), .QKV_weight_out_11_8(QKV_weight_out_11_8), .QKV_weight_out_11_9(QKV_weight_out_11_9), .QKV_weight_out_11_10(QKV_weight_out_11_10), .QKV_weight_out_11_11(QKV_weight_out_11_11), .QKV_weight_out_11_12(QKV_weight_out_11_12), .QKV_weight_out_11_13(QKV_weight_out_11_13), .QKV_weight_out_11_14(QKV_weight_out_11_14), .QKV_weight_out_11_15(QKV_weight_out_11_15),
    .QKV_weight_out_12_0(QKV_weight_out_12_0), .QKV_weight_out_12_1(QKV_weight_out_12_1), .QKV_weight_out_12_2(QKV_weight_out_12_2), .QKV_weight_out_12_3(QKV_weight_out_12_3), .QKV_weight_out_12_4(QKV_weight_out_12_4), .QKV_weight_out_12_5(QKV_weight_out_12_5), .QKV_weight_out_12_6(QKV_weight_out_12_6), .QKV_weight_out_12_7(QKV_weight_out_12_7), .QKV_weight_out_12_8(QKV_weight_out_12_8), .QKV_weight_out_12_9(QKV_weight_out_12_9), .QKV_weight_out_12_10(QKV_weight_out_12_10), .QKV_weight_out_12_11(QKV_weight_out_12_11), .QKV_weight_out_12_12(QKV_weight_out_12_12), .QKV_weight_out_12_13(QKV_weight_out_12_13), .QKV_weight_out_12_14(QKV_weight_out_12_14), .QKV_weight_out_12_15(QKV_weight_out_12_15),
    .QKV_weight_out_13_0(QKV_weight_out_13_0), .QKV_weight_out_13_1(QKV_weight_out_13_1), .QKV_weight_out_13_2(QKV_weight_out_13_2), .QKV_weight_out_13_3(QKV_weight_out_13_3), .QKV_weight_out_13_4(QKV_weight_out_13_4), .QKV_weight_out_13_5(QKV_weight_out_13_5), .QKV_weight_out_13_6(QKV_weight_out_13_6), .QKV_weight_out_13_7(QKV_weight_out_13_7), .QKV_weight_out_13_8(QKV_weight_out_13_8), .QKV_weight_out_13_9(QKV_weight_out_13_9), .QKV_weight_out_13_10(QKV_weight_out_13_10), .QKV_weight_out_13_11(QKV_weight_out_13_11), .QKV_weight_out_13_12(QKV_weight_out_13_12), .QKV_weight_out_13_13(QKV_weight_out_13_13), .QKV_weight_out_13_14(QKV_weight_out_13_14), .QKV_weight_out_13_15(QKV_weight_out_13_15),
    .QKV_weight_out_14_0(QKV_weight_out_14_0), .QKV_weight_out_14_1(QKV_weight_out_14_1), .QKV_weight_out_14_2(QKV_weight_out_14_2), .QKV_weight_out_14_3(QKV_weight_out_14_3), .QKV_weight_out_14_4(QKV_weight_out_14_4), .QKV_weight_out_14_5(QKV_weight_out_14_5), .QKV_weight_out_14_6(QKV_weight_out_14_6), .QKV_weight_out_14_7(QKV_weight_out_14_7), .QKV_weight_out_14_8(QKV_weight_out_14_8), .QKV_weight_out_14_9(QKV_weight_out_14_9), .QKV_weight_out_14_10(QKV_weight_out_14_10), .QKV_weight_out_14_11(QKV_weight_out_14_11), .QKV_weight_out_14_12(QKV_weight_out_14_12), .QKV_weight_out_14_13(QKV_weight_out_14_13), .QKV_weight_out_14_14(QKV_weight_out_14_14), .QKV_weight_out_14_15(QKV_weight_out_14_15),
    .QKV_weight_out_15_0(QKV_weight_out_15_0), .QKV_weight_out_15_1(QKV_weight_out_15_1), .QKV_weight_out_15_2(QKV_weight_out_15_2), .QKV_weight_out_15_3(QKV_weight_out_15_3), .QKV_weight_out_15_4(QKV_weight_out_15_4), .QKV_weight_out_15_5(QKV_weight_out_15_5), .QKV_weight_out_15_6(QKV_weight_out_15_6), .QKV_weight_out_15_7(QKV_weight_out_15_7), .QKV_weight_out_15_8(QKV_weight_out_15_8), .QKV_weight_out_15_9(QKV_weight_out_15_9), .QKV_weight_out_15_10(QKV_weight_out_15_10), .QKV_weight_out_15_11(QKV_weight_out_15_11), .QKV_weight_out_15_12(QKV_weight_out_15_12), .QKV_weight_out_15_13(QKV_weight_out_15_13), .QKV_weight_out_15_14(QKV_weight_out_15_14), .QKV_weight_out_15_15(QKV_weight_out_15_15),
    .QKV_weight_out_16_0(QKV_weight_out_16_0), .QKV_weight_out_16_1(QKV_weight_out_16_1), .QKV_weight_out_16_2(QKV_weight_out_16_2), .QKV_weight_out_16_3(QKV_weight_out_16_3), .QKV_weight_out_16_4(QKV_weight_out_16_4), .QKV_weight_out_16_5(QKV_weight_out_16_5), .QKV_weight_out_16_6(QKV_weight_out_16_6), .QKV_weight_out_16_7(QKV_weight_out_16_7), .QKV_weight_out_16_8(QKV_weight_out_16_8), .QKV_weight_out_16_9(QKV_weight_out_16_9), .QKV_weight_out_16_10(QKV_weight_out_16_10), .QKV_weight_out_16_11(QKV_weight_out_16_11), .QKV_weight_out_16_12(QKV_weight_out_16_12), .QKV_weight_out_16_13(QKV_weight_out_16_13), .QKV_weight_out_16_14(QKV_weight_out_16_14), .QKV_weight_out_16_15(QKV_weight_out_16_15),
    .QKV_weight_out_17_0(QKV_weight_out_17_0), .QKV_weight_out_17_1(QKV_weight_out_17_1), .QKV_weight_out_17_2(QKV_weight_out_17_2), .QKV_weight_out_17_3(QKV_weight_out_17_3), .QKV_weight_out_17_4(QKV_weight_out_17_4), .QKV_weight_out_17_5(QKV_weight_out_17_5), .QKV_weight_out_17_6(QKV_weight_out_17_6), .QKV_weight_out_17_7(QKV_weight_out_17_7), .QKV_weight_out_17_8(QKV_weight_out_17_8), .QKV_weight_out_17_9(QKV_weight_out_17_9), .QKV_weight_out_17_10(QKV_weight_out_17_10), .QKV_weight_out_17_11(QKV_weight_out_17_11), .QKV_weight_out_17_12(QKV_weight_out_17_12), .QKV_weight_out_17_13(QKV_weight_out_17_13), .QKV_weight_out_17_14(QKV_weight_out_17_14), .QKV_weight_out_17_15(QKV_weight_out_17_15),
    .QKV_weight_out_18_0(QKV_weight_out_18_0), .QKV_weight_out_18_1(QKV_weight_out_18_1), .QKV_weight_out_18_2(QKV_weight_out_18_2), .QKV_weight_out_18_3(QKV_weight_out_18_3), .QKV_weight_out_18_4(QKV_weight_out_18_4), .QKV_weight_out_18_5(QKV_weight_out_18_5), .QKV_weight_out_18_6(QKV_weight_out_18_6), .QKV_weight_out_18_7(QKV_weight_out_18_7), .QKV_weight_out_18_8(QKV_weight_out_18_8), .QKV_weight_out_18_9(QKV_weight_out_18_9), .QKV_weight_out_18_10(QKV_weight_out_18_10), .QKV_weight_out_18_11(QKV_weight_out_18_11), .QKV_weight_out_18_12(QKV_weight_out_18_12), .QKV_weight_out_18_13(QKV_weight_out_18_13), .QKV_weight_out_18_14(QKV_weight_out_18_14), .QKV_weight_out_18_15(QKV_weight_out_18_15),
    .QKV_weight_out_19_0(QKV_weight_out_19_0), .QKV_weight_out_19_1(QKV_weight_out_19_1), .QKV_weight_out_19_2(QKV_weight_out_19_2), .QKV_weight_out_19_3(QKV_weight_out_19_3), .QKV_weight_out_19_4(QKV_weight_out_19_4), .QKV_weight_out_19_5(QKV_weight_out_19_5), .QKV_weight_out_19_6(QKV_weight_out_19_6), .QKV_weight_out_19_7(QKV_weight_out_19_7), .QKV_weight_out_19_8(QKV_weight_out_19_8), .QKV_weight_out_19_9(QKV_weight_out_19_9), .QKV_weight_out_19_10(QKV_weight_out_19_10), .QKV_weight_out_19_11(QKV_weight_out_19_11), .QKV_weight_out_19_12(QKV_weight_out_19_12), .QKV_weight_out_19_13(QKV_weight_out_19_13), .QKV_weight_out_19_14(QKV_weight_out_19_14), .QKV_weight_out_19_15(QKV_weight_out_19_15),
    .QKV_weight_out_20_0(QKV_weight_out_20_0), .QKV_weight_out_20_1(QKV_weight_out_20_1), .QKV_weight_out_20_2(QKV_weight_out_20_2), .QKV_weight_out_20_3(QKV_weight_out_20_3), .QKV_weight_out_20_4(QKV_weight_out_20_4), .QKV_weight_out_20_5(QKV_weight_out_20_5), .QKV_weight_out_20_6(QKV_weight_out_20_6), .QKV_weight_out_20_7(QKV_weight_out_20_7), .QKV_weight_out_20_8(QKV_weight_out_20_8), .QKV_weight_out_20_9(QKV_weight_out_20_9), .QKV_weight_out_20_10(QKV_weight_out_20_10), .QKV_weight_out_20_11(QKV_weight_out_20_11), .QKV_weight_out_20_12(QKV_weight_out_20_12), .QKV_weight_out_20_13(QKV_weight_out_20_13), .QKV_weight_out_20_14(QKV_weight_out_20_14), .QKV_weight_out_20_15(QKV_weight_out_20_15),
    .QKV_weight_out_21_0(QKV_weight_out_21_0), .QKV_weight_out_21_1(QKV_weight_out_21_1), .QKV_weight_out_21_2(QKV_weight_out_21_2), .QKV_weight_out_21_3(QKV_weight_out_21_3), .QKV_weight_out_21_4(QKV_weight_out_21_4), .QKV_weight_out_21_5(QKV_weight_out_21_5), .QKV_weight_out_21_6(QKV_weight_out_21_6), .QKV_weight_out_21_7(QKV_weight_out_21_7), .QKV_weight_out_21_8(QKV_weight_out_21_8), .QKV_weight_out_21_9(QKV_weight_out_21_9), .QKV_weight_out_21_10(QKV_weight_out_21_10), .QKV_weight_out_21_11(QKV_weight_out_21_11), .QKV_weight_out_21_12(QKV_weight_out_21_12), .QKV_weight_out_21_13(QKV_weight_out_21_13), .QKV_weight_out_21_14(QKV_weight_out_21_14), .QKV_weight_out_21_15(QKV_weight_out_21_15),
    .QKV_weight_out_22_0(QKV_weight_out_22_0), .QKV_weight_out_22_1(QKV_weight_out_22_1), .QKV_weight_out_22_2(QKV_weight_out_22_2), .QKV_weight_out_22_3(QKV_weight_out_22_3), .QKV_weight_out_22_4(QKV_weight_out_22_4), .QKV_weight_out_22_5(QKV_weight_out_22_5), .QKV_weight_out_22_6(QKV_weight_out_22_6), .QKV_weight_out_22_7(QKV_weight_out_22_7), .QKV_weight_out_22_8(QKV_weight_out_22_8), .QKV_weight_out_22_9(QKV_weight_out_22_9), .QKV_weight_out_22_10(QKV_weight_out_22_10), .QKV_weight_out_22_11(QKV_weight_out_22_11), .QKV_weight_out_22_12(QKV_weight_out_22_12), .QKV_weight_out_22_13(QKV_weight_out_22_13), .QKV_weight_out_22_14(QKV_weight_out_22_14), .QKV_weight_out_22_15(QKV_weight_out_22_15),
    .QKV_weight_out_23_0(QKV_weight_out_23_0), .QKV_weight_out_23_1(QKV_weight_out_23_1), .QKV_weight_out_23_2(QKV_weight_out_23_2), .QKV_weight_out_23_3(QKV_weight_out_23_3), .QKV_weight_out_23_4(QKV_weight_out_23_4), .QKV_weight_out_23_5(QKV_weight_out_23_5), .QKV_weight_out_23_6(QKV_weight_out_23_6), .QKV_weight_out_23_7(QKV_weight_out_23_7), .QKV_weight_out_23_8(QKV_weight_out_23_8), .QKV_weight_out_23_9(QKV_weight_out_23_9), .QKV_weight_out_23_10(QKV_weight_out_23_10), .QKV_weight_out_23_11(QKV_weight_out_23_11), .QKV_weight_out_23_12(QKV_weight_out_23_12), .QKV_weight_out_23_13(QKV_weight_out_23_13), .QKV_weight_out_23_14(QKV_weight_out_23_14), .QKV_weight_out_23_15(QKV_weight_out_23_15),
    .QKV_weight_out_24_0(QKV_weight_out_24_0), .QKV_weight_out_24_1(QKV_weight_out_24_1), .QKV_weight_out_24_2(QKV_weight_out_24_2), .QKV_weight_out_24_3(QKV_weight_out_24_3), .QKV_weight_out_24_4(QKV_weight_out_24_4), .QKV_weight_out_24_5(QKV_weight_out_24_5), .QKV_weight_out_24_6(QKV_weight_out_24_6), .QKV_weight_out_24_7(QKV_weight_out_24_7), .QKV_weight_out_24_8(QKV_weight_out_24_8), .QKV_weight_out_24_9(QKV_weight_out_24_9), .QKV_weight_out_24_10(QKV_weight_out_24_10), .QKV_weight_out_24_11(QKV_weight_out_24_11), .QKV_weight_out_24_12(QKV_weight_out_24_12), .QKV_weight_out_24_13(QKV_weight_out_24_13), .QKV_weight_out_24_14(QKV_weight_out_24_14), .QKV_weight_out_24_15(QKV_weight_out_24_15),
    .QKV_weight_out_25_0(QKV_weight_out_25_0), .QKV_weight_out_25_1(QKV_weight_out_25_1), .QKV_weight_out_25_2(QKV_weight_out_25_2), .QKV_weight_out_25_3(QKV_weight_out_25_3), .QKV_weight_out_25_4(QKV_weight_out_25_4), .QKV_weight_out_25_5(QKV_weight_out_25_5), .QKV_weight_out_25_6(QKV_weight_out_25_6), .QKV_weight_out_25_7(QKV_weight_out_25_7), .QKV_weight_out_25_8(QKV_weight_out_25_8), .QKV_weight_out_25_9(QKV_weight_out_25_9), .QKV_weight_out_25_10(QKV_weight_out_25_10), .QKV_weight_out_25_11(QKV_weight_out_25_11), .QKV_weight_out_25_12(QKV_weight_out_25_12), .QKV_weight_out_25_13(QKV_weight_out_25_13), .QKV_weight_out_25_14(QKV_weight_out_25_14), .QKV_weight_out_25_15(QKV_weight_out_25_15),
    .QKV_weight_out_26_0(QKV_weight_out_26_0), .QKV_weight_out_26_1(QKV_weight_out_26_1), .QKV_weight_out_26_2(QKV_weight_out_26_2), .QKV_weight_out_26_3(QKV_weight_out_26_3), .QKV_weight_out_26_4(QKV_weight_out_26_4), .QKV_weight_out_26_5(QKV_weight_out_26_5), .QKV_weight_out_26_6(QKV_weight_out_26_6), .QKV_weight_out_26_7(QKV_weight_out_26_7), .QKV_weight_out_26_8(QKV_weight_out_26_8), .QKV_weight_out_26_9(QKV_weight_out_26_9), .QKV_weight_out_26_10(QKV_weight_out_26_10), .QKV_weight_out_26_11(QKV_weight_out_26_11), .QKV_weight_out_26_12(QKV_weight_out_26_12), .QKV_weight_out_26_13(QKV_weight_out_26_13), .QKV_weight_out_26_14(QKV_weight_out_26_14), .QKV_weight_out_26_15(QKV_weight_out_26_15),
    .QKV_weight_out_27_0(QKV_weight_out_27_0), .QKV_weight_out_27_1(QKV_weight_out_27_1), .QKV_weight_out_27_2(QKV_weight_out_27_2), .QKV_weight_out_27_3(QKV_weight_out_27_3), .QKV_weight_out_27_4(QKV_weight_out_27_4), .QKV_weight_out_27_5(QKV_weight_out_27_5), .QKV_weight_out_27_6(QKV_weight_out_27_6), .QKV_weight_out_27_7(QKV_weight_out_27_7), .QKV_weight_out_27_8(QKV_weight_out_27_8), .QKV_weight_out_27_9(QKV_weight_out_27_9), .QKV_weight_out_27_10(QKV_weight_out_27_10), .QKV_weight_out_27_11(QKV_weight_out_27_11), .QKV_weight_out_27_12(QKV_weight_out_27_12), .QKV_weight_out_27_13(QKV_weight_out_27_13), .QKV_weight_out_27_14(QKV_weight_out_27_14), .QKV_weight_out_27_15(QKV_weight_out_27_15),
    .QKV_weight_out_28_0(QKV_weight_out_28_0), .QKV_weight_out_28_1(QKV_weight_out_28_1), .QKV_weight_out_28_2(QKV_weight_out_28_2), .QKV_weight_out_28_3(QKV_weight_out_28_3), .QKV_weight_out_28_4(QKV_weight_out_28_4), .QKV_weight_out_28_5(QKV_weight_out_28_5), .QKV_weight_out_28_6(QKV_weight_out_28_6), .QKV_weight_out_28_7(QKV_weight_out_28_7), .QKV_weight_out_28_8(QKV_weight_out_28_8), .QKV_weight_out_28_9(QKV_weight_out_28_9), .QKV_weight_out_28_10(QKV_weight_out_28_10), .QKV_weight_out_28_11(QKV_weight_out_28_11), .QKV_weight_out_28_12(QKV_weight_out_28_12), .QKV_weight_out_28_13(QKV_weight_out_28_13), .QKV_weight_out_28_14(QKV_weight_out_28_14), .QKV_weight_out_28_15(QKV_weight_out_28_15),
    .QKV_weight_out_29_0(QKV_weight_out_29_0), .QKV_weight_out_29_1(QKV_weight_out_29_1), .QKV_weight_out_29_2(QKV_weight_out_29_2), .QKV_weight_out_29_3(QKV_weight_out_29_3), .QKV_weight_out_29_4(QKV_weight_out_29_4), .QKV_weight_out_29_5(QKV_weight_out_29_5), .QKV_weight_out_29_6(QKV_weight_out_29_6), .QKV_weight_out_29_7(QKV_weight_out_29_7), .QKV_weight_out_29_8(QKV_weight_out_29_8), .QKV_weight_out_29_9(QKV_weight_out_29_9), .QKV_weight_out_29_10(QKV_weight_out_29_10), .QKV_weight_out_29_11(QKV_weight_out_29_11), .QKV_weight_out_29_12(QKV_weight_out_29_12), .QKV_weight_out_29_13(QKV_weight_out_29_13), .QKV_weight_out_29_14(QKV_weight_out_29_14), .QKV_weight_out_29_15(QKV_weight_out_29_15),
    .QKV_weight_out_30_0(QKV_weight_out_30_0), .QKV_weight_out_30_1(QKV_weight_out_30_1), .QKV_weight_out_30_2(QKV_weight_out_30_2), .QKV_weight_out_30_3(QKV_weight_out_30_3), .QKV_weight_out_30_4(QKV_weight_out_30_4), .QKV_weight_out_30_5(QKV_weight_out_30_5), .QKV_weight_out_30_6(QKV_weight_out_30_6), .QKV_weight_out_30_7(QKV_weight_out_30_7), .QKV_weight_out_30_8(QKV_weight_out_30_8), .QKV_weight_out_30_9(QKV_weight_out_30_9), .QKV_weight_out_30_10(QKV_weight_out_30_10), .QKV_weight_out_30_11(QKV_weight_out_30_11), .QKV_weight_out_30_12(QKV_weight_out_30_12), .QKV_weight_out_30_13(QKV_weight_out_30_13), .QKV_weight_out_30_14(QKV_weight_out_30_14), .QKV_weight_out_30_15(QKV_weight_out_30_15),
    .QKV_weight_out_31_0(QKV_weight_out_31_0), .QKV_weight_out_31_1(QKV_weight_out_31_1), .QKV_weight_out_31_2(QKV_weight_out_31_2), .QKV_weight_out_31_3(QKV_weight_out_31_3), .QKV_weight_out_31_4(QKV_weight_out_31_4), .QKV_weight_out_31_5(QKV_weight_out_31_5), .QKV_weight_out_31_6(QKV_weight_out_31_6), .QKV_weight_out_31_7(QKV_weight_out_31_7), .QKV_weight_out_31_8(QKV_weight_out_31_8), .QKV_weight_out_31_9(QKV_weight_out_31_9), .QKV_weight_out_31_10(QKV_weight_out_31_10), .QKV_weight_out_31_11(QKV_weight_out_31_11), .QKV_weight_out_31_12(QKV_weight_out_31_12), .QKV_weight_out_31_13(QKV_weight_out_31_13), .QKV_weight_out_31_14(QKV_weight_out_31_14), .QKV_weight_out_31_15(QKV_weight_out_31_15),
    
    .QKT_weight_out_0_0(QKT_weight_out_0_0), .QKT_weight_out_0_1(QKT_weight_out_0_1), .QKT_weight_out_0_2(QKT_weight_out_0_2), .QKT_weight_out_0_3(QKT_weight_out_0_3), .QKT_weight_out_0_4(QKT_weight_out_0_4), .QKT_weight_out_0_5(QKT_weight_out_0_5), .QKT_weight_out_0_6(QKT_weight_out_0_6), .QKT_weight_out_0_7(QKT_weight_out_0_7), .QKT_weight_out_0_8(QKT_weight_out_0_8), .QKT_weight_out_0_9(QKT_weight_out_0_9), .QKT_weight_out_0_10(QKT_weight_out_0_10), .QKT_weight_out_0_11(QKT_weight_out_0_11), .QKT_weight_out_0_12(QKT_weight_out_0_12), .QKT_weight_out_0_13(QKT_weight_out_0_13), .QKT_weight_out_0_14(QKT_weight_out_0_14), .QKT_weight_out_0_15(QKT_weight_out_0_15),
    .QKT_weight_out_1_0(QKT_weight_out_1_0), .QKT_weight_out_1_1(QKT_weight_out_1_1), .QKT_weight_out_1_2(QKT_weight_out_1_2), .QKT_weight_out_1_3(QKT_weight_out_1_3), .QKT_weight_out_1_4(QKT_weight_out_1_4), .QKT_weight_out_1_5(QKT_weight_out_1_5), .QKT_weight_out_1_6(QKT_weight_out_1_6), .QKT_weight_out_1_7(QKT_weight_out_1_7), .QKT_weight_out_1_8(QKT_weight_out_1_8), .QKT_weight_out_1_9(QKT_weight_out_1_9), .QKT_weight_out_1_10(QKT_weight_out_1_10), .QKT_weight_out_1_11(QKT_weight_out_1_11), .QKT_weight_out_1_12(QKT_weight_out_1_12), .QKT_weight_out_1_13(QKT_weight_out_1_13), .QKT_weight_out_1_14(QKT_weight_out_1_14), .QKT_weight_out_1_15(QKT_weight_out_1_15),
    .QKT_weight_out_2_0(QKT_weight_out_2_0), .QKT_weight_out_2_1(QKT_weight_out_2_1), .QKT_weight_out_2_2(QKT_weight_out_2_2), .QKT_weight_out_2_3(QKT_weight_out_2_3), .QKT_weight_out_2_4(QKT_weight_out_2_4), .QKT_weight_out_2_5(QKT_weight_out_2_5), .QKT_weight_out_2_6(QKT_weight_out_2_6), .QKT_weight_out_2_7(QKT_weight_out_2_7), .QKT_weight_out_2_8(QKT_weight_out_2_8), .QKT_weight_out_2_9(QKT_weight_out_2_9), .QKT_weight_out_2_10(QKT_weight_out_2_10), .QKT_weight_out_2_11(QKT_weight_out_2_11), .QKT_weight_out_2_12(QKT_weight_out_2_12), .QKT_weight_out_2_13(QKT_weight_out_2_13), .QKT_weight_out_2_14(QKT_weight_out_2_14), .QKT_weight_out_2_15(QKT_weight_out_2_15),
    .QKT_weight_out_3_0(QKT_weight_out_3_0), .QKT_weight_out_3_1(QKT_weight_out_3_1), .QKT_weight_out_3_2(QKT_weight_out_3_2), .QKT_weight_out_3_3(QKT_weight_out_3_3), .QKT_weight_out_3_4(QKT_weight_out_3_4), .QKT_weight_out_3_5(QKT_weight_out_3_5), .QKT_weight_out_3_6(QKT_weight_out_3_6), .QKT_weight_out_3_7(QKT_weight_out_3_7), .QKT_weight_out_3_8(QKT_weight_out_3_8), .QKT_weight_out_3_9(QKT_weight_out_3_9), .QKT_weight_out_3_10(QKT_weight_out_3_10), .QKT_weight_out_3_11(QKT_weight_out_3_11), .QKT_weight_out_3_12(QKT_weight_out_3_12), .QKT_weight_out_3_13(QKT_weight_out_3_13), .QKT_weight_out_3_14(QKT_weight_out_3_14), .QKT_weight_out_3_15(QKT_weight_out_3_15),

    .QKV_data_out_0_0(QKV_data_out_0_0), .QKV_data_out_0_1(QKV_data_out_0_1), .QKV_data_out_0_2(QKV_data_out_0_2), .QKV_data_out_0_3(QKV_data_out_0_3), .QKV_data_out_0_4(QKV_data_out_0_4), .QKV_data_out_0_5(QKV_data_out_0_5), .QKV_data_out_0_6(QKV_data_out_0_6), .QKV_data_out_0_7(QKV_data_out_0_7), .QKV_data_out_0_8(QKV_data_out_0_8), .QKV_data_out_0_9(QKV_data_out_0_9), .QKV_data_out_0_10(QKV_data_out_0_10), .QKV_data_out_0_11(QKV_data_out_0_11), .QKV_data_out_0_12(QKV_data_out_0_12), .QKV_data_out_0_13(QKV_data_out_0_13), .QKV_data_out_0_14(QKV_data_out_0_14), .QKV_data_out_0_15(QKV_data_out_0_15),
    .QKV_data_out_1_0(QKV_data_out_1_0), .QKV_data_out_1_1(QKV_data_out_1_1), .QKV_data_out_1_2(QKV_data_out_1_2), .QKV_data_out_1_3(QKV_data_out_1_3), .QKV_data_out_1_4(QKV_data_out_1_4), .QKV_data_out_1_5(QKV_data_out_1_5), .QKV_data_out_1_6(QKV_data_out_1_6), .QKV_data_out_1_7(QKV_data_out_1_7), .QKV_data_out_1_8(QKV_data_out_1_8), .QKV_data_out_1_9(QKV_data_out_1_9), .QKV_data_out_1_10(QKV_data_out_1_10), .QKV_data_out_1_11(QKV_data_out_1_11), .QKV_data_out_1_12(QKV_data_out_1_12), .QKV_data_out_1_13(QKV_data_out_1_13), .QKV_data_out_1_14(QKV_data_out_1_14), .QKV_data_out_1_15(QKV_data_out_1_15),
    .QKV_data_out_2_0(QKV_data_out_2_0), .QKV_data_out_2_1(QKV_data_out_2_1), .QKV_data_out_2_2(QKV_data_out_2_2), .QKV_data_out_2_3(QKV_data_out_2_3), .QKV_data_out_2_4(QKV_data_out_2_4), .QKV_data_out_2_5(QKV_data_out_2_5), .QKV_data_out_2_6(QKV_data_out_2_6), .QKV_data_out_2_7(QKV_data_out_2_7), .QKV_data_out_2_8(QKV_data_out_2_8), .QKV_data_out_2_9(QKV_data_out_2_9), .QKV_data_out_2_10(QKV_data_out_2_10), .QKV_data_out_2_11(QKV_data_out_2_11), .QKV_data_out_2_12(QKV_data_out_2_12), .QKV_data_out_2_13(QKV_data_out_2_13), .QKV_data_out_2_14(QKV_data_out_2_14), .QKV_data_out_2_15(QKV_data_out_2_15),
    .QKV_data_out_3_0(QKV_data_out_3_0), .QKV_data_out_3_1(QKV_data_out_3_1), .QKV_data_out_3_2(QKV_data_out_3_2), .QKV_data_out_3_3(QKV_data_out_3_3), .QKV_data_out_3_4(QKV_data_out_3_4), .QKV_data_out_3_5(QKV_data_out_3_5), .QKV_data_out_3_6(QKV_data_out_3_6), .QKV_data_out_3_7(QKV_data_out_3_7), .QKV_data_out_3_8(QKV_data_out_3_8), .QKV_data_out_3_9(QKV_data_out_3_9), .QKV_data_out_3_10(QKV_data_out_3_10), .QKV_data_out_3_11(QKV_data_out_3_11), .QKV_data_out_3_12(QKV_data_out_3_12), .QKV_data_out_3_13(QKV_data_out_3_13), .QKV_data_out_3_14(QKV_data_out_3_14), .QKV_data_out_3_15(QKV_data_out_3_15),
    .QKV_data_out_4_0(QKV_data_out_4_0), .QKV_data_out_4_1(QKV_data_out_4_1), .QKV_data_out_4_2(QKV_data_out_4_2), .QKV_data_out_4_3(QKV_data_out_4_3), .QKV_data_out_4_4(QKV_data_out_4_4), .QKV_data_out_4_5(QKV_data_out_4_5), .QKV_data_out_4_6(QKV_data_out_4_6), .QKV_data_out_4_7(QKV_data_out_4_7), .QKV_data_out_4_8(QKV_data_out_4_8), .QKV_data_out_4_9(QKV_data_out_4_9), .QKV_data_out_4_10(QKV_data_out_4_10), .QKV_data_out_4_11(QKV_data_out_4_11), .QKV_data_out_4_12(QKV_data_out_4_12), .QKV_data_out_4_13(QKV_data_out_4_13), .QKV_data_out_4_14(QKV_data_out_4_14), .QKV_data_out_4_15(QKV_data_out_4_15),
    .QKV_data_out_5_0(QKV_data_out_5_0), .QKV_data_out_5_1(QKV_data_out_5_1), .QKV_data_out_5_2(QKV_data_out_5_2), .QKV_data_out_5_3(QKV_data_out_5_3), .QKV_data_out_5_4(QKV_data_out_5_4), .QKV_data_out_5_5(QKV_data_out_5_5), .QKV_data_out_5_6(QKV_data_out_5_6), .QKV_data_out_5_7(QKV_data_out_5_7), .QKV_data_out_5_8(QKV_data_out_5_8), .QKV_data_out_5_9(QKV_data_out_5_9), .QKV_data_out_5_10(QKV_data_out_5_10), .QKV_data_out_5_11(QKV_data_out_5_11), .QKV_data_out_5_12(QKV_data_out_5_12), .QKV_data_out_5_13(QKV_data_out_5_13), .QKV_data_out_5_14(QKV_data_out_5_14), .QKV_data_out_5_15(QKV_data_out_5_15),
    .QKV_data_out_6_0(QKV_data_out_6_0), .QKV_data_out_6_1(QKV_data_out_6_1), .QKV_data_out_6_2(QKV_data_out_6_2), .QKV_data_out_6_3(QKV_data_out_6_3), .QKV_data_out_6_4(QKV_data_out_6_4), .QKV_data_out_6_5(QKV_data_out_6_5), .QKV_data_out_6_6(QKV_data_out_6_6), .QKV_data_out_6_7(QKV_data_out_6_7), .QKV_data_out_6_8(QKV_data_out_6_8), .QKV_data_out_6_9(QKV_data_out_6_9), .QKV_data_out_6_10(QKV_data_out_6_10), .QKV_data_out_6_11(QKV_data_out_6_11), .QKV_data_out_6_12(QKV_data_out_6_12), .QKV_data_out_6_13(QKV_data_out_6_13), .QKV_data_out_6_14(QKV_data_out_6_14), .QKV_data_out_6_15(QKV_data_out_6_15),
    .QKV_data_out_7_0(QKV_data_out_7_0), .QKV_data_out_7_1(QKV_data_out_7_1), .QKV_data_out_7_2(QKV_data_out_7_2), .QKV_data_out_7_3(QKV_data_out_7_3), .QKV_data_out_7_4(QKV_data_out_7_4), .QKV_data_out_7_5(QKV_data_out_7_5), .QKV_data_out_7_6(QKV_data_out_7_6), .QKV_data_out_7_7(QKV_data_out_7_7), .QKV_data_out_7_8(QKV_data_out_7_8), .QKV_data_out_7_9(QKV_data_out_7_9), .QKV_data_out_7_10(QKV_data_out_7_10), .QKV_data_out_7_11(QKV_data_out_7_11), .QKV_data_out_7_12(QKV_data_out_7_12), .QKV_data_out_7_13(QKV_data_out_7_13), .QKV_data_out_7_14(QKV_data_out_7_14), .QKV_data_out_7_15(QKV_data_out_7_15),
    .QKV_data_out_8_0(QKV_data_out_8_0), .QKV_data_out_8_1(QKV_data_out_8_1), .QKV_data_out_8_2(QKV_data_out_8_2), .QKV_data_out_8_3(QKV_data_out_8_3), .QKV_data_out_8_4(QKV_data_out_8_4), .QKV_data_out_8_5(QKV_data_out_8_5), .QKV_data_out_8_6(QKV_data_out_8_6), .QKV_data_out_8_7(QKV_data_out_8_7), .QKV_data_out_8_8(QKV_data_out_8_8), .QKV_data_out_8_9(QKV_data_out_8_9), .QKV_data_out_8_10(QKV_data_out_8_10), .QKV_data_out_8_11(QKV_data_out_8_11), .QKV_data_out_8_12(QKV_data_out_8_12), .QKV_data_out_8_13(QKV_data_out_8_13), .QKV_data_out_8_14(QKV_data_out_8_14), .QKV_data_out_8_15(QKV_data_out_8_15),
    .QKV_data_out_9_0(QKV_data_out_9_0), .QKV_data_out_9_1(QKV_data_out_9_1), .QKV_data_out_9_2(QKV_data_out_9_2), .QKV_data_out_9_3(QKV_data_out_9_3), .QKV_data_out_9_4(QKV_data_out_9_4), .QKV_data_out_9_5(QKV_data_out_9_5), .QKV_data_out_9_6(QKV_data_out_9_6), .QKV_data_out_9_7(QKV_data_out_9_7), .QKV_data_out_9_8(QKV_data_out_9_8), .QKV_data_out_9_9(QKV_data_out_9_9), .QKV_data_out_9_10(QKV_data_out_9_10), .QKV_data_out_9_11(QKV_data_out_9_11), .QKV_data_out_9_12(QKV_data_out_9_12), .QKV_data_out_9_13(QKV_data_out_9_13), .QKV_data_out_9_14(QKV_data_out_9_14), .QKV_data_out_9_15(QKV_data_out_9_15),
    .QKV_data_out_10_0(QKV_data_out_10_0), .QKV_data_out_10_1(QKV_data_out_10_1), .QKV_data_out_10_2(QKV_data_out_10_2), .QKV_data_out_10_3(QKV_data_out_10_3), .QKV_data_out_10_4(QKV_data_out_10_4), .QKV_data_out_10_5(QKV_data_out_10_5), .QKV_data_out_10_6(QKV_data_out_10_6), .QKV_data_out_10_7(QKV_data_out_10_7), .QKV_data_out_10_8(QKV_data_out_10_8), .QKV_data_out_10_9(QKV_data_out_10_9), .QKV_data_out_10_10(QKV_data_out_10_10), .QKV_data_out_10_11(QKV_data_out_10_11), .QKV_data_out_10_12(QKV_data_out_10_12), .QKV_data_out_10_13(QKV_data_out_10_13), .QKV_data_out_10_14(QKV_data_out_10_14), .QKV_data_out_10_15(QKV_data_out_10_15),
    .QKV_data_out_11_0(QKV_data_out_11_0), .QKV_data_out_11_1(QKV_data_out_11_1), .QKV_data_out_11_2(QKV_data_out_11_2), .QKV_data_out_11_3(QKV_data_out_11_3), .QKV_data_out_11_4(QKV_data_out_11_4), .QKV_data_out_11_5(QKV_data_out_11_5), .QKV_data_out_11_6(QKV_data_out_11_6), .QKV_data_out_11_7(QKV_data_out_11_7), .QKV_data_out_11_8(QKV_data_out_11_8), .QKV_data_out_11_9(QKV_data_out_11_9), .QKV_data_out_11_10(QKV_data_out_11_10), .QKV_data_out_11_11(QKV_data_out_11_11), .QKV_data_out_11_12(QKV_data_out_11_12), .QKV_data_out_11_13(QKV_data_out_11_13), .QKV_data_out_11_14(QKV_data_out_11_14), .QKV_data_out_11_15(QKV_data_out_11_15),
    .QKV_data_out_12_0(QKV_data_out_12_0), .QKV_data_out_12_1(QKV_data_out_12_1), .QKV_data_out_12_2(QKV_data_out_12_2), .QKV_data_out_12_3(QKV_data_out_12_3), .QKV_data_out_12_4(QKV_data_out_12_4), .QKV_data_out_12_5(QKV_data_out_12_5), .QKV_data_out_12_6(QKV_data_out_12_6), .QKV_data_out_12_7(QKV_data_out_12_7), .QKV_data_out_12_8(QKV_data_out_12_8), .QKV_data_out_12_9(QKV_data_out_12_9), .QKV_data_out_12_10(QKV_data_out_12_10), .QKV_data_out_12_11(QKV_data_out_12_11), .QKV_data_out_12_12(QKV_data_out_12_12), .QKV_data_out_12_13(QKV_data_out_12_13), .QKV_data_out_12_14(QKV_data_out_12_14), .QKV_data_out_12_15(QKV_data_out_12_15),
    .QKV_data_out_13_0(QKV_data_out_13_0), .QKV_data_out_13_1(QKV_data_out_13_1), .QKV_data_out_13_2(QKV_data_out_13_2), .QKV_data_out_13_3(QKV_data_out_13_3), .QKV_data_out_13_4(QKV_data_out_13_4), .QKV_data_out_13_5(QKV_data_out_13_5), .QKV_data_out_13_6(QKV_data_out_13_6), .QKV_data_out_13_7(QKV_data_out_13_7), .QKV_data_out_13_8(QKV_data_out_13_8), .QKV_data_out_13_9(QKV_data_out_13_9), .QKV_data_out_13_10(QKV_data_out_13_10), .QKV_data_out_13_11(QKV_data_out_13_11), .QKV_data_out_13_12(QKV_data_out_13_12), .QKV_data_out_13_13(QKV_data_out_13_13), .QKV_data_out_13_14(QKV_data_out_13_14), .QKV_data_out_13_15(QKV_data_out_13_15),
    .QKV_data_out_14_0(QKV_data_out_14_0), .QKV_data_out_14_1(QKV_data_out_14_1), .QKV_data_out_14_2(QKV_data_out_14_2), .QKV_data_out_14_3(QKV_data_out_14_3), .QKV_data_out_14_4(QKV_data_out_14_4), .QKV_data_out_14_5(QKV_data_out_14_5), .QKV_data_out_14_6(QKV_data_out_14_6), .QKV_data_out_14_7(QKV_data_out_14_7), .QKV_data_out_14_8(QKV_data_out_14_8), .QKV_data_out_14_9(QKV_data_out_14_9), .QKV_data_out_14_10(QKV_data_out_14_10), .QKV_data_out_14_11(QKV_data_out_14_11), .QKV_data_out_14_12(QKV_data_out_14_12), .QKV_data_out_14_13(QKV_data_out_14_13), .QKV_data_out_14_14(QKV_data_out_14_14), .QKV_data_out_14_15(QKV_data_out_14_15),
    .QKV_data_out_15_0(QKV_data_out_15_0), .QKV_data_out_15_1(QKV_data_out_15_1), .QKV_data_out_15_2(QKV_data_out_15_2), .QKV_data_out_15_3(QKV_data_out_15_3), .QKV_data_out_15_4(QKV_data_out_15_4), .QKV_data_out_15_5(QKV_data_out_15_5), .QKV_data_out_15_6(QKV_data_out_15_6), .QKV_data_out_15_7(QKV_data_out_15_7), .QKV_data_out_15_8(QKV_data_out_15_8), .QKV_data_out_15_9(QKV_data_out_15_9), .QKV_data_out_15_10(QKV_data_out_15_10), .QKV_data_out_15_11(QKV_data_out_15_11), .QKV_data_out_15_12(QKV_data_out_15_12), .QKV_data_out_15_13(QKV_data_out_15_13), .QKV_data_out_15_14(QKV_data_out_15_14), .QKV_data_out_15_15(QKV_data_out_15_15),
    .QKV_data_out_16_0(QKV_data_out_16_0), .QKV_data_out_16_1(QKV_data_out_16_1), .QKV_data_out_16_2(QKV_data_out_16_2), .QKV_data_out_16_3(QKV_data_out_16_3), .QKV_data_out_16_4(QKV_data_out_16_4), .QKV_data_out_16_5(QKV_data_out_16_5), .QKV_data_out_16_6(QKV_data_out_16_6), .QKV_data_out_16_7(QKV_data_out_16_7), .QKV_data_out_16_8(QKV_data_out_16_8), .QKV_data_out_16_9(QKV_data_out_16_9), .QKV_data_out_16_10(QKV_data_out_16_10), .QKV_data_out_16_11(QKV_data_out_16_11), .QKV_data_out_16_12(QKV_data_out_16_12), .QKV_data_out_16_13(QKV_data_out_16_13), .QKV_data_out_16_14(QKV_data_out_16_14), .QKV_data_out_16_15(QKV_data_out_16_15),
    .QKV_data_out_17_0(QKV_data_out_17_0), .QKV_data_out_17_1(QKV_data_out_17_1), .QKV_data_out_17_2(QKV_data_out_17_2), .QKV_data_out_17_3(QKV_data_out_17_3), .QKV_data_out_17_4(QKV_data_out_17_4), .QKV_data_out_17_5(QKV_data_out_17_5), .QKV_data_out_17_6(QKV_data_out_17_6), .QKV_data_out_17_7(QKV_data_out_17_7), .QKV_data_out_17_8(QKV_data_out_17_8), .QKV_data_out_17_9(QKV_data_out_17_9), .QKV_data_out_17_10(QKV_data_out_17_10), .QKV_data_out_17_11(QKV_data_out_17_11), .QKV_data_out_17_12(QKV_data_out_17_12), .QKV_data_out_17_13(QKV_data_out_17_13), .QKV_data_out_17_14(QKV_data_out_17_14), .QKV_data_out_17_15(QKV_data_out_17_15),
    .QKV_data_out_18_0(QKV_data_out_18_0), .QKV_data_out_18_1(QKV_data_out_18_1), .QKV_data_out_18_2(QKV_data_out_18_2), .QKV_data_out_18_3(QKV_data_out_18_3), .QKV_data_out_18_4(QKV_data_out_18_4), .QKV_data_out_18_5(QKV_data_out_18_5), .QKV_data_out_18_6(QKV_data_out_18_6), .QKV_data_out_18_7(QKV_data_out_18_7), .QKV_data_out_18_8(QKV_data_out_18_8), .QKV_data_out_18_9(QKV_data_out_18_9), .QKV_data_out_18_10(QKV_data_out_18_10), .QKV_data_out_18_11(QKV_data_out_18_11), .QKV_data_out_18_12(QKV_data_out_18_12), .QKV_data_out_18_13(QKV_data_out_18_13), .QKV_data_out_18_14(QKV_data_out_18_14), .QKV_data_out_18_15(QKV_data_out_18_15),
    .QKV_data_out_19_0(QKV_data_out_19_0), .QKV_data_out_19_1(QKV_data_out_19_1), .QKV_data_out_19_2(QKV_data_out_19_2), .QKV_data_out_19_3(QKV_data_out_19_3), .QKV_data_out_19_4(QKV_data_out_19_4), .QKV_data_out_19_5(QKV_data_out_19_5), .QKV_data_out_19_6(QKV_data_out_19_6), .QKV_data_out_19_7(QKV_data_out_19_7), .QKV_data_out_19_8(QKV_data_out_19_8), .QKV_data_out_19_9(QKV_data_out_19_9), .QKV_data_out_19_10(QKV_data_out_19_10), .QKV_data_out_19_11(QKV_data_out_19_11), .QKV_data_out_19_12(QKV_data_out_19_12), .QKV_data_out_19_13(QKV_data_out_19_13), .QKV_data_out_19_14(QKV_data_out_19_14), .QKV_data_out_19_15(QKV_data_out_19_15),
    .QKV_data_out_20_0(QKV_data_out_20_0), .QKV_data_out_20_1(QKV_data_out_20_1), .QKV_data_out_20_2(QKV_data_out_20_2), .QKV_data_out_20_3(QKV_data_out_20_3), .QKV_data_out_20_4(QKV_data_out_20_4), .QKV_data_out_20_5(QKV_data_out_20_5), .QKV_data_out_20_6(QKV_data_out_20_6), .QKV_data_out_20_7(QKV_data_out_20_7), .QKV_data_out_20_8(QKV_data_out_20_8), .QKV_data_out_20_9(QKV_data_out_20_9), .QKV_data_out_20_10(QKV_data_out_20_10), .QKV_data_out_20_11(QKV_data_out_20_11), .QKV_data_out_20_12(QKV_data_out_20_12), .QKV_data_out_20_13(QKV_data_out_20_13), .QKV_data_out_20_14(QKV_data_out_20_14), .QKV_data_out_20_15(QKV_data_out_20_15),
    .QKV_data_out_21_0(QKV_data_out_21_0), .QKV_data_out_21_1(QKV_data_out_21_1), .QKV_data_out_21_2(QKV_data_out_21_2), .QKV_data_out_21_3(QKV_data_out_21_3), .QKV_data_out_21_4(QKV_data_out_21_4), .QKV_data_out_21_5(QKV_data_out_21_5), .QKV_data_out_21_6(QKV_data_out_21_6), .QKV_data_out_21_7(QKV_data_out_21_7), .QKV_data_out_21_8(QKV_data_out_21_8), .QKV_data_out_21_9(QKV_data_out_21_9), .QKV_data_out_21_10(QKV_data_out_21_10), .QKV_data_out_21_11(QKV_data_out_21_11), .QKV_data_out_21_12(QKV_data_out_21_12), .QKV_data_out_21_13(QKV_data_out_21_13), .QKV_data_out_21_14(QKV_data_out_21_14), .QKV_data_out_21_15(QKV_data_out_21_15),
    .QKV_data_out_22_0(QKV_data_out_22_0), .QKV_data_out_22_1(QKV_data_out_22_1), .QKV_data_out_22_2(QKV_data_out_22_2), .QKV_data_out_22_3(QKV_data_out_22_3), .QKV_data_out_22_4(QKV_data_out_22_4), .QKV_data_out_22_5(QKV_data_out_22_5), .QKV_data_out_22_6(QKV_data_out_22_6), .QKV_data_out_22_7(QKV_data_out_22_7), .QKV_data_out_22_8(QKV_data_out_22_8), .QKV_data_out_22_9(QKV_data_out_22_9), .QKV_data_out_22_10(QKV_data_out_22_10), .QKV_data_out_22_11(QKV_data_out_22_11), .QKV_data_out_22_12(QKV_data_out_22_12), .QKV_data_out_22_13(QKV_data_out_22_13), .QKV_data_out_22_14(QKV_data_out_22_14), .QKV_data_out_22_15(QKV_data_out_22_15),
    .QKV_data_out_23_0(QKV_data_out_23_0), .QKV_data_out_23_1(QKV_data_out_23_1), .QKV_data_out_23_2(QKV_data_out_23_2), .QKV_data_out_23_3(QKV_data_out_23_3), .QKV_data_out_23_4(QKV_data_out_23_4), .QKV_data_out_23_5(QKV_data_out_23_5), .QKV_data_out_23_6(QKV_data_out_23_6), .QKV_data_out_23_7(QKV_data_out_23_7), .QKV_data_out_23_8(QKV_data_out_23_8), .QKV_data_out_23_9(QKV_data_out_23_9), .QKV_data_out_23_10(QKV_data_out_23_10), .QKV_data_out_23_11(QKV_data_out_23_11), .QKV_data_out_23_12(QKV_data_out_23_12), .QKV_data_out_23_13(QKV_data_out_23_13), .QKV_data_out_23_14(QKV_data_out_23_14), .QKV_data_out_23_15(QKV_data_out_23_15),
    .QKV_data_out_24_0(QKV_data_out_24_0), .QKV_data_out_24_1(QKV_data_out_24_1), .QKV_data_out_24_2(QKV_data_out_24_2), .QKV_data_out_24_3(QKV_data_out_24_3), .QKV_data_out_24_4(QKV_data_out_24_4), .QKV_data_out_24_5(QKV_data_out_24_5), .QKV_data_out_24_6(QKV_data_out_24_6), .QKV_data_out_24_7(QKV_data_out_24_7), .QKV_data_out_24_8(QKV_data_out_24_8), .QKV_data_out_24_9(QKV_data_out_24_9), .QKV_data_out_24_10(QKV_data_out_24_10), .QKV_data_out_24_11(QKV_data_out_24_11), .QKV_data_out_24_12(QKV_data_out_24_12), .QKV_data_out_24_13(QKV_data_out_24_13), .QKV_data_out_24_14(QKV_data_out_24_14), .QKV_data_out_24_15(QKV_data_out_24_15),
    .QKV_data_out_25_0(QKV_data_out_25_0), .QKV_data_out_25_1(QKV_data_out_25_1), .QKV_data_out_25_2(QKV_data_out_25_2), .QKV_data_out_25_3(QKV_data_out_25_3), .QKV_data_out_25_4(QKV_data_out_25_4), .QKV_data_out_25_5(QKV_data_out_25_5), .QKV_data_out_25_6(QKV_data_out_25_6), .QKV_data_out_25_7(QKV_data_out_25_7), .QKV_data_out_25_8(QKV_data_out_25_8), .QKV_data_out_25_9(QKV_data_out_25_9), .QKV_data_out_25_10(QKV_data_out_25_10), .QKV_data_out_25_11(QKV_data_out_25_11), .QKV_data_out_25_12(QKV_data_out_25_12), .QKV_data_out_25_13(QKV_data_out_25_13), .QKV_data_out_25_14(QKV_data_out_25_14), .QKV_data_out_25_15(QKV_data_out_25_15),
    .QKV_data_out_26_0(QKV_data_out_26_0), .QKV_data_out_26_1(QKV_data_out_26_1), .QKV_data_out_26_2(QKV_data_out_26_2), .QKV_data_out_26_3(QKV_data_out_26_3), .QKV_data_out_26_4(QKV_data_out_26_4), .QKV_data_out_26_5(QKV_data_out_26_5), .QKV_data_out_26_6(QKV_data_out_26_6), .QKV_data_out_26_7(QKV_data_out_26_7), .QKV_data_out_26_8(QKV_data_out_26_8), .QKV_data_out_26_9(QKV_data_out_26_9), .QKV_data_out_26_10(QKV_data_out_26_10), .QKV_data_out_26_11(QKV_data_out_26_11), .QKV_data_out_26_12(QKV_data_out_26_12), .QKV_data_out_26_13(QKV_data_out_26_13), .QKV_data_out_26_14(QKV_data_out_26_14), .QKV_data_out_26_15(QKV_data_out_26_15),
    .QKV_data_out_27_0(QKV_data_out_27_0), .QKV_data_out_27_1(QKV_data_out_27_1), .QKV_data_out_27_2(QKV_data_out_27_2), .QKV_data_out_27_3(QKV_data_out_27_3), .QKV_data_out_27_4(QKV_data_out_27_4), .QKV_data_out_27_5(QKV_data_out_27_5), .QKV_data_out_27_6(QKV_data_out_27_6), .QKV_data_out_27_7(QKV_data_out_27_7), .QKV_data_out_27_8(QKV_data_out_27_8), .QKV_data_out_27_9(QKV_data_out_27_9), .QKV_data_out_27_10(QKV_data_out_27_10), .QKV_data_out_27_11(QKV_data_out_27_11), .QKV_data_out_27_12(QKV_data_out_27_12), .QKV_data_out_27_13(QKV_data_out_27_13), .QKV_data_out_27_14(QKV_data_out_27_14), .QKV_data_out_27_15(QKV_data_out_27_15),
    .QKV_data_out_28_0(QKV_data_out_28_0), .QKV_data_out_28_1(QKV_data_out_28_1), .QKV_data_out_28_2(QKV_data_out_28_2), .QKV_data_out_28_3(QKV_data_out_28_3), .QKV_data_out_28_4(QKV_data_out_28_4), .QKV_data_out_28_5(QKV_data_out_28_5), .QKV_data_out_28_6(QKV_data_out_28_6), .QKV_data_out_28_7(QKV_data_out_28_7), .QKV_data_out_28_8(QKV_data_out_28_8), .QKV_data_out_28_9(QKV_data_out_28_9), .QKV_data_out_28_10(QKV_data_out_28_10), .QKV_data_out_28_11(QKV_data_out_28_11), .QKV_data_out_28_12(QKV_data_out_28_12), .QKV_data_out_28_13(QKV_data_out_28_13), .QKV_data_out_28_14(QKV_data_out_28_14), .QKV_data_out_28_15(QKV_data_out_28_15),
    .QKV_data_out_29_0(QKV_data_out_29_0), .QKV_data_out_29_1(QKV_data_out_29_1), .QKV_data_out_29_2(QKV_data_out_29_2), .QKV_data_out_29_3(QKV_data_out_29_3), .QKV_data_out_29_4(QKV_data_out_29_4), .QKV_data_out_29_5(QKV_data_out_29_5), .QKV_data_out_29_6(QKV_data_out_29_6), .QKV_data_out_29_7(QKV_data_out_29_7), .QKV_data_out_29_8(QKV_data_out_29_8), .QKV_data_out_29_9(QKV_data_out_29_9), .QKV_data_out_29_10(QKV_data_out_29_10), .QKV_data_out_29_11(QKV_data_out_29_11), .QKV_data_out_29_12(QKV_data_out_29_12), .QKV_data_out_29_13(QKV_data_out_29_13), .QKV_data_out_29_14(QKV_data_out_29_14), .QKV_data_out_29_15(QKV_data_out_29_15),
    .QKV_data_out_30_0(QKV_data_out_30_0), .QKV_data_out_30_1(QKV_data_out_30_1), .QKV_data_out_30_2(QKV_data_out_30_2), .QKV_data_out_30_3(QKV_data_out_30_3), .QKV_data_out_30_4(QKV_data_out_30_4), .QKV_data_out_30_5(QKV_data_out_30_5), .QKV_data_out_30_6(QKV_data_out_30_6), .QKV_data_out_30_7(QKV_data_out_30_7), .QKV_data_out_30_8(QKV_data_out_30_8), .QKV_data_out_30_9(QKV_data_out_30_9), .QKV_data_out_30_10(QKV_data_out_30_10), .QKV_data_out_30_11(QKV_data_out_30_11), .QKV_data_out_30_12(QKV_data_out_30_12), .QKV_data_out_30_13(QKV_data_out_30_13), .QKV_data_out_30_14(QKV_data_out_30_14), .QKV_data_out_30_15(QKV_data_out_30_15),
    .QKV_data_out_31_0(QKV_data_out_31_0), .QKV_data_out_31_1(QKV_data_out_31_1), .QKV_data_out_31_2(QKV_data_out_31_2), .QKV_data_out_31_3(QKV_data_out_31_3), .QKV_data_out_31_4(QKV_data_out_31_4), .QKV_data_out_31_5(QKV_data_out_31_5), .QKV_data_out_31_6(QKV_data_out_31_6), .QKV_data_out_31_7(QKV_data_out_31_7), .QKV_data_out_31_8(QKV_data_out_31_8), .QKV_data_out_31_9(QKV_data_out_31_9), .QKV_data_out_31_10(QKV_data_out_31_10), .QKV_data_out_31_11(QKV_data_out_31_11), .QKV_data_out_31_12(QKV_data_out_31_12), .QKV_data_out_31_13(QKV_data_out_31_13), .QKV_data_out_31_14(QKV_data_out_31_14), .QKV_data_out_31_15(QKV_data_out_31_15),

    .QKT_data_out_0_0(QKT_data_out_0_0), .QKT_data_out_0_1(QKT_data_out_0_1), .QKT_data_out_0_2(QKT_data_out_0_2), .QKT_data_out_0_3(QKT_data_out_0_3), .QKT_data_out_0_4(QKT_data_out_0_4), .QKT_data_out_0_5(QKT_data_out_0_5), .QKT_data_out_0_6(QKT_data_out_0_6), .QKT_data_out_0_7(QKT_data_out_0_7), .QKT_data_out_0_8(QKT_data_out_0_8), .QKT_data_out_0_9(QKT_data_out_0_9), .QKT_data_out_0_10(QKT_data_out_0_10), .QKT_data_out_0_11(QKT_data_out_0_11), .QKT_data_out_0_12(QKT_data_out_0_12), .QKT_data_out_0_13(QKT_data_out_0_13), .QKT_data_out_0_14(QKT_data_out_0_14), .QKT_data_out_0_15(QKT_data_out_0_15),
    .QKT_data_out_1_0(QKT_data_out_1_0), .QKT_data_out_1_1(QKT_data_out_1_1), .QKT_data_out_1_2(QKT_data_out_1_2), .QKT_data_out_1_3(QKT_data_out_1_3), .QKT_data_out_1_4(QKT_data_out_1_4), .QKT_data_out_1_5(QKT_data_out_1_5), .QKT_data_out_1_6(QKT_data_out_1_6), .QKT_data_out_1_7(QKT_data_out_1_7), .QKT_data_out_1_8(QKT_data_out_1_8), .QKT_data_out_1_9(QKT_data_out_1_9), .QKT_data_out_1_10(QKT_data_out_1_10), .QKT_data_out_1_11(QKT_data_out_1_11), .QKT_data_out_1_12(QKT_data_out_1_12), .QKT_data_out_1_13(QKT_data_out_1_13), .QKT_data_out_1_14(QKT_data_out_1_14), .QKT_data_out_1_15(QKT_data_out_1_15),
    .QKT_data_out_2_0(QKT_data_out_2_0), .QKT_data_out_2_1(QKT_data_out_2_1), .QKT_data_out_2_2(QKT_data_out_2_2), .QKT_data_out_2_3(QKT_data_out_2_3), .QKT_data_out_2_4(QKT_data_out_2_4), .QKT_data_out_2_5(QKT_data_out_2_5), .QKT_data_out_2_6(QKT_data_out_2_6), .QKT_data_out_2_7(QKT_data_out_2_7), .QKT_data_out_2_8(QKT_data_out_2_8), .QKT_data_out_2_9(QKT_data_out_2_9), .QKT_data_out_2_10(QKT_data_out_2_10), .QKT_data_out_2_11(QKT_data_out_2_11), .QKT_data_out_2_12(QKT_data_out_2_12), .QKT_data_out_2_13(QKT_data_out_2_13), .QKT_data_out_2_14(QKT_data_out_2_14), .QKT_data_out_2_15(QKT_data_out_2_15),
    .QKT_data_out_3_0(QKT_data_out_3_0), .QKT_data_out_3_1(QKT_data_out_3_1), .QKT_data_out_3_2(QKT_data_out_3_2), .QKT_data_out_3_3(QKT_data_out_3_3), .QKT_data_out_3_4(QKT_data_out_3_4), .QKT_data_out_3_5(QKT_data_out_3_5), .QKT_data_out_3_6(QKT_data_out_3_6), .QKT_data_out_3_7(QKT_data_out_3_7), .QKT_data_out_3_8(QKT_data_out_3_8), .QKT_data_out_3_9(QKT_data_out_3_9), .QKT_data_out_3_10(QKT_data_out_3_10), .QKT_data_out_3_11(QKT_data_out_3_11), .QKT_data_out_3_12(QKT_data_out_3_12), .QKT_data_out_3_13(QKT_data_out_3_13), .QKT_data_out_3_14(QKT_data_out_3_14), .QKT_data_out_3_15(QKT_data_out_3_15),

    .QKV_is_write_out_0(QKV_is_write_out_0), .QKV_is_write_out_1(QKV_is_write_out_1), .QKV_is_write_out_2(QKV_is_write_out_2), .QKV_is_write_out_3(QKV_is_write_out_3), .QKV_is_write_out_4(QKV_is_write_out_4), .QKV_is_write_out_5(QKV_is_write_out_5), .QKV_is_write_out_6(QKV_is_write_out_6), .QKV_is_write_out_7(QKV_is_write_out_7), .QKV_is_write_out_8(QKV_is_write_out_8), .QKV_is_write_out_9(QKV_is_write_out_9), .QKV_is_write_out_10(QKV_is_write_out_10), .QKV_is_write_out_11(QKV_is_write_out_11), .QKV_is_write_out_12(QKV_is_write_out_12), .QKV_is_write_out_13(QKV_is_write_out_13), .QKV_is_write_out_14(QKV_is_write_out_14), 
    .QKV_is_write_out_15(QKV_is_write_out_15), .QKV_is_write_out_16(QKV_is_write_out_16), .QKV_is_write_out_17(QKV_is_write_out_17), .QKV_is_write_out_18(QKV_is_write_out_18), .QKV_is_write_out_19(QKV_is_write_out_19), .QKV_is_write_out_20(QKV_is_write_out_20), .QKV_is_write_out_21(QKV_is_write_out_21), .QKV_is_write_out_22(QKV_is_write_out_22), .QKV_is_write_out_23(QKV_is_write_out_23), .QKV_is_write_out_24(QKV_is_write_out_24), .QKV_is_write_out_25(QKV_is_write_out_25), .QKV_is_write_out_26(QKV_is_write_out_26), .QKV_is_write_out_27(QKV_is_write_out_27), .QKV_is_write_out_28(QKV_is_write_out_28), .QKV_is_write_out_29(QKV_is_write_out_29), .QKV_is_write_out_30(QKV_is_write_out_30), .QKV_is_write_out_31(QKV_is_write_out_31), 

    .QKV_selcet_out_0(QKV_selcet_out_0), .QKV_selcet_out_1(QKV_selcet_out_1), .QKV_selcet_out_2(QKV_selcet_out_2), .QKV_selcet_out_3(QKV_selcet_out_3), .QKV_selcet_out_4(QKV_selcet_out_4), .QKV_selcet_out_5(QKV_selcet_out_5), .QKV_selcet_out_6(QKV_selcet_out_6), .QKV_selcet_out_7(QKV_selcet_out_7), .QKV_selcet_out_8(QKV_selcet_out_8), .QKV_selcet_out_9(QKV_selcet_out_9), .QKV_selcet_out_10(QKV_selcet_out_10), .QKV_selcet_out_11(QKV_selcet_out_11), .QKV_selcet_out_12(QKV_selcet_out_12), .QKV_selcet_out_13(QKV_selcet_out_13), .QKV_selcet_out_14(QKV_selcet_out_14), .QKV_selcet_out_15(QKV_selcet_out_15), 
    .QKV_selcet_out_16(QKV_selcet_out_16), .QKV_selcet_out_17(QKV_selcet_out_17), .QKV_selcet_out_18(QKV_selcet_out_18), .QKV_selcet_out_19(QKV_selcet_out_19), .QKV_selcet_out_20(QKV_selcet_out_20), .QKV_selcet_out_21(QKV_selcet_out_21), .QKV_selcet_out_22(QKV_selcet_out_22), .QKV_selcet_out_23(QKV_selcet_out_23), .QKV_selcet_out_24(QKV_selcet_out_24), .QKV_selcet_out_25(QKV_selcet_out_25), .QKV_selcet_out_26(QKV_selcet_out_26), .QKV_selcet_out_27(QKV_selcet_out_27), .QKV_selcet_out_28(QKV_selcet_out_28), .QKV_selcet_out_29(QKV_selcet_out_29), .QKV_selcet_out_30(QKV_selcet_out_30), .QKV_selcet_out_31(QKV_selcet_out_31),

    .QKT_is_write_out_0(QKT_is_write_out_0), .QKT_is_write_out_1(QKT_is_write_out_1), .QKT_is_write_out_2(QKT_is_write_out_2), .QKT_is_write_out_3(QKT_is_write_out_3), 

    .QKT_select_out_0(QKT_select_out_0), .QKT_select_out_1(QKT_select_out_1), .QKT_select_out_2(QKT_select_out_2), .QKT_select_out_3(QKT_select_out_3), 


);

dimc_macro i_dimc_macro_0(.input_addr(QKV_addr_out_0), 
                          .input_weight_0(QKV_weight_out_0_0), .input_weight_1(QKV_weight_out_0_1), .input_weight_2(QKV_weight_out_0_2), .input_weight_3(QKV_weight_out_0_3), .input_weight_4(QKV_weight_out_0_4), .input_weight_5(QKV_weight_out_0_5), .input_weight_6(QKV_weight_out_0_6), .input_weight_7(QKV_weight_out_0_7), .input_weight_8(QKV_weight_out_0_8), .input_weight_9(QKV_weight_out_0_9), .input_weight_10(QKV_weight_out_0_10), .input_weight_11(QKV_weight_out_0_11), .input_weight_12(QKV_weight_out_0_12), .input_weight_13(QKV_weight_out_0_13), .input_weight_14(QKV_weight_out_0_14), .input_weight_15(QKV_weight_out_0_15),
                          .input_data_0(QKV_data_out_0_0), .input_data_1(QKV_data_out_0_1), .input_data_2(QKV_data_out_0_2), .input_data_3(QKV_data_out_0_3), .input_data_4(QKV_data_out_0_4), .input_data_5(QKV_data_out_0_5), .input_data_6(QKV_data_out_0_6), .input_data_7(QKV_data_out_0_7), .input_data_8(QKV_data_out_0_8), .input_data_9(QKV_data_out_0_9), .input_data_10(QKV_data_out_0_10), .input_data_11(QKV_data_out_0_11), .input_data_12(QKV_data_out_0_12), .input_data_13(QKV_data_out_0_13), .input_data_14(QKV_data_out_0_14), .input_data_15(QKV_data_out_0_15),
                          .is_write_(QKV_is_write_out_0), .select_(QKV_selcet_out_0),
                          .calc_result_0(QKV_calc_result_0_0), .calc_result_1(QKV_calc_result_0_1), .calc_result_2(QKV_calc_result_0_2), .calc_result_3(QKV_calc_result_0_3), .calc_result_4(QKV_calc_result_0_4), .calc_result_5(QKV_calc_result_0_5), .calc_result_6(QKV_calc_result_0_6), .calc_result_7(QKV_calc_result_0_7), .calc_result_8(QKV_calc_result_0_8), .calc_result_9(QKV_calc_result_0_9), .calc_result_10(QKV_calc_result_0_10), .calc_result_11(QKV_calc_result_0_11), .calc_result_12(QKV_calc_result_0_12), .calc_result_13(QKV_calc_result_0_13), .calc_result_14(QKV_calc_result_0_14), .calc_result_15(QKV_calc_result_0_15)
);

dimc_macro i_dimc_macro_0(.input_addr(QKV_addr_out_0),
                          .input_weight_0(QKV_weight_out_0_0), .input_weight_1(QKV_weight_out_0_1), .input_weight_2(QKV_weight_out_0_2), .input_weight_3(QKV_weight_out_0_3), .input_weight_4(QKV_weight_out_0_4), .input_weight_5(QKV_weight_out_0_5), .input_weight_6(QKV_weight_out_0_6), .input_weight_7(QKV_weight_out_0_7), .input_weight_8(QKV_weight_out_0_8), .input_weight_9(QKV_weight_out_0_9), .input_weight_10(QKV_weight_out_0_10), .input_weight_11(QKV_weight_out_0_11), .input_weight_12(QKV_weight_out_0_12), .input_weight_13(QKV_weight_out_0_13), .input_weight_14(QKV_weight_out_0_14), .input_weight_15(QKV_weight_out_0_15),
                          .input_data_0(QKV_data_out_0_0), .input_data_1(QKV_data_out_0_1), .input_data_2(QKV_data_out_0_2), .input_data_3(QKV_data_out_0_3), .input_data_4(QKV_data_out_0_4), .input_data_5(QKV_data_out_0_5), .input_data_6(QKV_data_out_0_6), .input_data_7(QKV_data_out_0_7), .input_data_8(QKV_data_out_0_8), .input_data_9(QKV_data_out_0_9), .input_data_10(QKV_data_out_0_10), .input_data_11(QKV_data_out_0_11), .input_data_12(QKV_data_out_0_12), .input_data_13(QKV_data_out_0_13), .input_data_14(QKV_data_out_0_14), .input_data_15(QKV_data_out_0_15),
                          .is_write_(QKV_is_write_out_0), .select_(QKV_selcet_out_0),
                          .calc_result_0(QKV_calc_result_0_0), .calc_result_1(QKV_calc_result_0_1), .calc_result_2(QKV_calc_result_0_2), .calc_result_3(QKV_calc_result_0_3), .calc_result_4(QKV_calc_result_0_4), .calc_result_5(QKV_calc_result_0_5), .calc_result_6(QKV_calc_result_0_6), .calc_result_7(QKV_calc_result_0_7), .calc_result_8(QKV_calc_result_0_8), .calc_result_9(QKV_calc_result_0_9), .calc_result_10(QKV_calc_result_0_10), .calc_result_11(QKV_calc_result_0_11), .calc_result_12(QKV_calc_result_0_12), .calc_result_13(QKV_calc_result_0_13), .calc_result_14(QKV_calc_result_0_14), .calc_result_15(QKV_calc_result_0_15)
);

dimc_macro i_dimc_macro_1(.input_addr(QKV_addr_out_1),
                          .input_weight_0(QKV_weight_out_1_0), .input_weight_1(QKV_weight_out_1_1), .input_weight_2(QKV_weight_out_1_2), .input_weight_3(QKV_weight_out_1_3), .input_weight_4(QKV_weight_out_1_4), .input_weight_5(QKV_weight_out_1_5), .input_weight_6(QKV_weight_out_1_6), .input_weight_7(QKV_weight_out_1_7), .input_weight_8(QKV_weight_out_1_8), .input_weight_9(QKV_weight_out_1_9), .input_weight_10(QKV_weight_out_1_10), .input_weight_11(QKV_weight_out_1_11), .input_weight_12(QKV_weight_out_1_12), .input_weight_13(QKV_weight_out_1_13), .input_weight_14(QKV_weight_out_1_14), .input_weight_15(QKV_weight_out_1_15),
                          .input_data_0(QKV_data_out_1_0), .input_data_1(QKV_data_out_1_1), .input_data_2(QKV_data_out_1_2), .input_data_3(QKV_data_out_1_3), .input_data_4(QKV_data_out_1_4), .input_data_5(QKV_data_out_1_5), .input_data_6(QKV_data_out_1_6), .input_data_7(QKV_data_out_1_7), .input_data_8(QKV_data_out_1_8), .input_data_9(QKV_data_out_1_9), .input_data_10(QKV_data_out_1_10), .input_data_11(QKV_data_out_1_11), .input_data_12(QKV_data_out_1_12), .input_data_13(QKV_data_out_1_13), .input_data_14(QKV_data_out_1_14), .input_data_15(QKV_data_out_1_15),
                          .is_write_(QKV_is_write_out_1), .select_(QKV_selcet_out_1),
                          .calc_result_0(QKV_calc_result_1_0), .calc_result_1(QKV_calc_result_1_1), .calc_result_2(QKV_calc_result_1_2), .calc_result_3(QKV_calc_result_1_3), .calc_result_4(QKV_calc_result_1_4), .calc_result_5(QKV_calc_result_1_5), .calc_result_6(QKV_calc_result_1_6), .calc_result_7(QKV_calc_result_1_7), .calc_result_8(QKV_calc_result_1_8), .calc_result_9(QKV_calc_result_1_9), .calc_result_10(QKV_calc_result_1_10), .calc_result_11(QKV_calc_result_1_11), .calc_result_12(QKV_calc_result_1_12), .calc_result_13(QKV_calc_result_1_13), .calc_result_14(QKV_calc_result_1_14), .calc_result_15(QKV_calc_result_1_15)
);

dimc_macro i_dimc_macro_2(.input_addr(QKV_addr_out_2),
                          .input_weight_0(QKV_weight_out_2_0), .input_weight_1(QKV_weight_out_2_1), .input_weight_2(QKV_weight_out_2_2), .input_weight_3(QKV_weight_out_2_3), .input_weight_4(QKV_weight_out_2_4), .input_weight_5(QKV_weight_out_2_5), .input_weight_6(QKV_weight_out_2_6), .input_weight_7(QKV_weight_out_2_7), .input_weight_8(QKV_weight_out_2_8), .input_weight_9(QKV_weight_out_2_9), .input_weight_10(QKV_weight_out_2_10), .input_weight_11(QKV_weight_out_2_11), .input_weight_12(QKV_weight_out_2_12), .input_weight_13(QKV_weight_out_2_13), .input_weight_14(QKV_weight_out_2_14), .input_weight_15(QKV_weight_out_2_15),
                          .input_data_0(QKV_data_out_2_0), .input_data_1(QKV_data_out_2_1), .input_data_2(QKV_data_out_2_2), .input_data_3(QKV_data_out_2_3), .input_data_4(QKV_data_out_2_4), .input_data_5(QKV_data_out_2_5), .input_data_6(QKV_data_out_2_6), .input_data_7(QKV_data_out_2_7), .input_data_8(QKV_data_out_2_8), .input_data_9(QKV_data_out_2_9), .input_data_10(QKV_data_out_2_10), .input_data_11(QKV_data_out_2_11), .input_data_12(QKV_data_out_2_12), .input_data_13(QKV_data_out_2_13), .input_data_14(QKV_data_out_2_14), .input_data_15(QKV_data_out_2_15),
                          .is_write_(QKV_is_write_out_2), .select_(QKV_selcet_out_2),
                          .calc_result_0(QKV_calc_result_2_0), .calc_result_1(QKV_calc_result_2_1), .calc_result_2(QKV_calc_result_2_2), .calc_result_3(QKV_calc_result_2_3), .calc_result_4(QKV_calc_result_2_4), .calc_result_5(QKV_calc_result_2_5), .calc_result_6(QKV_calc_result_2_6), .calc_result_7(QKV_calc_result_2_7), .calc_result_8(QKV_calc_result_2_8), .calc_result_9(QKV_calc_result_2_9), .calc_result_10(QKV_calc_result_2_10), .calc_result_11(QKV_calc_result_2_11), .calc_result_12(QKV_calc_result_2_12), .calc_result_13(QKV_calc_result_2_13), .calc_result_14(QKV_calc_result_2_14), .calc_result_15(QKV_calc_result_2_15)
);

dimc_macro i_dimc_macro_3(.input_addr(QKV_addr_out_3),
                          .input_weight_0(QKV_weight_out_3_0), .input_weight_1(QKV_weight_out_3_1), .input_weight_2(QKV_weight_out_3_2), .input_weight_3(QKV_weight_out_3_3), .input_weight_4(QKV_weight_out_3_4), .input_weight_5(QKV_weight_out_3_5), .input_weight_6(QKV_weight_out_3_6), .input_weight_7(QKV_weight_out_3_7), .input_weight_8(QKV_weight_out_3_8), .input_weight_9(QKV_weight_out_3_9), .input_weight_10(QKV_weight_out_3_10), .input_weight_11(QKV_weight_out_3_11), .input_weight_12(QKV_weight_out_3_12), .input_weight_13(QKV_weight_out_3_13), .input_weight_14(QKV_weight_out_3_14), .input_weight_15(QKV_weight_out_3_15),
                          .input_data_0(QKV_data_out_3_0), .input_data_1(QKV_data_out_3_1), .input_data_2(QKV_data_out_3_2), .input_data_3(QKV_data_out_3_3), .input_data_4(QKV_data_out_3_4), .input_data_5(QKV_data_out_3_5), .input_data_6(QKV_data_out_3_6), .input_data_7(QKV_data_out_3_7), .input_data_8(QKV_data_out_3_8), .input_data_9(QKV_data_out_3_9), .input_data_10(QKV_data_out_3_10), .input_data_11(QKV_data_out_3_11), .input_data_12(QKV_data_out_3_12), .input_data_13(QKV_data_out_3_13), .input_data_14(QKV_data_out_3_14), .input_data_15(QKV_data_out_3_15),
                          .is_write_(QKV_is_write_out_3), .select_(QKV_selcet_out_3),
                          .calc_result_0(QKV_calc_result_3_0), .calc_result_1(QKV_calc_result_3_1), .calc_result_2(QKV_calc_result_3_2), .calc_result_3(QKV_calc_result_3_3), .calc_result_4(QKV_calc_result_3_4), .calc_result_5(QKV_calc_result_3_5), .calc_result_6(QKV_calc_result_3_6), .calc_result_7(QKV_calc_result_3_7), .calc_result_8(QKV_calc_result_3_8), .calc_result_9(QKV_calc_result_3_9), .calc_result_10(QKV_calc_result_3_10), .calc_result_11(QKV_calc_result_3_11), .calc_result_12(QKV_calc_result_3_12), .calc_result_13(QKV_calc_result_3_13), .calc_result_14(QKV_calc_result_3_14), .calc_result_15(QKV_calc_result_3_15)
);

dimc_macro i_dimc_macro_4(.input_addr(QKV_addr_out_4),
                          .input_weight_0(QKV_weight_out_4_0), .input_weight_1(QKV_weight_out_4_1), .input_weight_2(QKV_weight_out_4_2), .input_weight_3(QKV_weight_out_4_3), .input_weight_4(QKV_weight_out_4_4), .input_weight_5(QKV_weight_out_4_5), .input_weight_6(QKV_weight_out_4_6), .input_weight_7(QKV_weight_out_4_7), .input_weight_8(QKV_weight_out_4_8), .input_weight_9(QKV_weight_out_4_9), .input_weight_10(QKV_weight_out_4_10), .input_weight_11(QKV_weight_out_4_11), .input_weight_12(QKV_weight_out_4_12), .input_weight_13(QKV_weight_out_4_13), .input_weight_14(QKV_weight_out_4_14), .input_weight_15(QKV_weight_out_4_15),
                          .input_data_0(QKV_data_out_4_0), .input_data_1(QKV_data_out_4_1), .input_data_2(QKV_data_out_4_2), .input_data_3(QKV_data_out_4_3), .input_data_4(QKV_data_out_4_4), .input_data_5(QKV_data_out_4_5), .input_data_6(QKV_data_out_4_6), .input_data_7(QKV_data_out_4_7), .input_data_8(QKV_data_out_4_8), .input_data_9(QKV_data_out_4_9), .input_data_10(QKV_data_out_4_10), .input_data_11(QKV_data_out_4_11), .input_data_12(QKV_data_out_4_12), .input_data_13(QKV_data_out_4_13), .input_data_14(QKV_data_out_4_14), .input_data_15(QKV_data_out_4_15),
                          .is_write_(QKV_is_write_out_4), .select_(QKV_selcet_out_4),
                          .calc_result_0(QKV_calc_result_4_0), .calc_result_1(QKV_calc_result_4_1), .calc_result_2(QKV_calc_result_4_2), .calc_result_3(QKV_calc_result_4_3), .calc_result_4(QKV_calc_result_4_4), .calc_result_5(QKV_calc_result_4_5), .calc_result_6(QKV_calc_result_4_6), .calc_result_7(QKV_calc_result_4_7), .calc_result_8(QKV_calc_result_4_8), .calc_result_9(QKV_calc_result_4_9), .calc_result_10(QKV_calc_result_4_10), .calc_result_11(QKV_calc_result_4_11), .calc_result_12(QKV_calc_result_4_12), .calc_result_13(QKV_calc_result_4_13), .calc_result_14(QKV_calc_result_4_14), .calc_result_15(QKV_calc_result_4_15)
);

dimc_macro i_dimc_macro_5(.input_addr(QKV_addr_out_5),
                          .input_weight_0(QKV_weight_out_5_0), .input_weight_1(QKV_weight_out_5_1), .input_weight_2(QKV_weight_out_5_2), .input_weight_3(QKV_weight_out_5_3), .input_weight_4(QKV_weight_out_5_4), .input_weight_5(QKV_weight_out_5_5), .input_weight_6(QKV_weight_out_5_6), .input_weight_7(QKV_weight_out_5_7), .input_weight_8(QKV_weight_out_5_8), .input_weight_9(QKV_weight_out_5_9), .input_weight_10(QKV_weight_out_5_10), .input_weight_11(QKV_weight_out_5_11), .input_weight_12(QKV_weight_out_5_12), .input_weight_13(QKV_weight_out_5_13), .input_weight_14(QKV_weight_out_5_14), .input_weight_15(QKV_weight_out_5_15),
                          .input_data_0(QKV_data_out_5_0), .input_data_1(QKV_data_out_5_1), .input_data_2(QKV_data_out_5_2), .input_data_3(QKV_data_out_5_3), .input_data_4(QKV_data_out_5_4), .input_data_5(QKV_data_out_5_5), .input_data_6(QKV_data_out_5_6), .input_data_7(QKV_data_out_5_7), .input_data_8(QKV_data_out_5_8), .input_data_9(QKV_data_out_5_9), .input_data_10(QKV_data_out_5_10), .input_data_11(QKV_data_out_5_11), .input_data_12(QKV_data_out_5_12), .input_data_13(QKV_data_out_5_13), .input_data_14(QKV_data_out_5_14), .input_data_15(QKV_data_out_5_15),
                          .is_write_(QKV_is_write_out_5), .select_(QKV_selcet_out_5),
                          .calc_result_0(QKV_calc_result_5_0), .calc_result_1(QKV_calc_result_5_1), .calc_result_2(QKV_calc_result_5_2), .calc_result_3(QKV_calc_result_5_3), .calc_result_4(QKV_calc_result_5_4), .calc_result_5(QKV_calc_result_5_5), .calc_result_6(QKV_calc_result_5_6), .calc_result_7(QKV_calc_result_5_7), .calc_result_8(QKV_calc_result_5_8), .calc_result_9(QKV_calc_result_5_9), .calc_result_10(QKV_calc_result_5_10), .calc_result_11(QKV_calc_result_5_11), .calc_result_12(QKV_calc_result_5_12), .calc_result_13(QKV_calc_result_5_13), .calc_result_14(QKV_calc_result_5_14), .calc_result_15(QKV_calc_result_5_15)
);

dimc_macro i_dimc_macro_6(.input_addr(QKV_addr_out_6),
                          .input_weight_0(QKV_weight_out_6_0), .input_weight_1(QKV_weight_out_6_1), .input_weight_2(QKV_weight_out_6_2), .input_weight_3(QKV_weight_out_6_3), .input_weight_4(QKV_weight_out_6_4), .input_weight_5(QKV_weight_out_6_5), .input_weight_6(QKV_weight_out_6_6), .input_weight_7(QKV_weight_out_6_7), .input_weight_8(QKV_weight_out_6_8), .input_weight_9(QKV_weight_out_6_9), .input_weight_10(QKV_weight_out_6_10), .input_weight_11(QKV_weight_out_6_11), .input_weight_12(QKV_weight_out_6_12), .input_weight_13(QKV_weight_out_6_13), .input_weight_14(QKV_weight_out_6_14), .input_weight_15(QKV_weight_out_6_15),
                          .input_data_0(QKV_data_out_6_0), .input_data_1(QKV_data_out_6_1), .input_data_2(QKV_data_out_6_2), .input_data_3(QKV_data_out_6_3), .input_data_4(QKV_data_out_6_4), .input_data_5(QKV_data_out_6_5), .input_data_6(QKV_data_out_6_6), .input_data_7(QKV_data_out_6_7), .input_data_8(QKV_data_out_6_8), .input_data_9(QKV_data_out_6_9), .input_data_10(QKV_data_out_6_10), .input_data_11(QKV_data_out_6_11), .input_data_12(QKV_data_out_6_12), .input_data_13(QKV_data_out_6_13), .input_data_14(QKV_data_out_6_14), .input_data_15(QKV_data_out_6_15),
                          .is_write_(QKV_is_write_out_6), .select_(QKV_selcet_out_6),
                          .calc_result_0(QKV_calc_result_6_0), .calc_result_1(QKV_calc_result_6_1), .calc_result_2(QKV_calc_result_6_2), .calc_result_3(QKV_calc_result_6_3), .calc_result_4(QKV_calc_result_6_4), .calc_result_5(QKV_calc_result_6_5), .calc_result_6(QKV_calc_result_6_6), .calc_result_7(QKV_calc_result_6_7), .calc_result_8(QKV_calc_result_6_8), .calc_result_9(QKV_calc_result_6_9), .calc_result_10(QKV_calc_result_6_10), .calc_result_11(QKV_calc_result_6_11), .calc_result_12(QKV_calc_result_6_12), .calc_result_13(QKV_calc_result_6_13), .calc_result_14(QKV_calc_result_6_14), .calc_result_15(QKV_calc_result_6_15)
);

dimc_macro i_dimc_macro_7(.input_addr(QKV_addr_out_7),
                          .input_weight_0(QKV_weight_out_7_0), .input_weight_1(QKV_weight_out_7_1), .input_weight_2(QKV_weight_out_7_2), .input_weight_3(QKV_weight_out_7_3), .input_weight_4(QKV_weight_out_7_4), .input_weight_5(QKV_weight_out_7_5), .input_weight_6(QKV_weight_out_7_6), .input_weight_7(QKV_weight_out_7_7), .input_weight_8(QKV_weight_out_7_8), .input_weight_9(QKV_weight_out_7_9), .input_weight_10(QKV_weight_out_7_10), .input_weight_11(QKV_weight_out_7_11), .input_weight_12(QKV_weight_out_7_12), .input_weight_13(QKV_weight_out_7_13), .input_weight_14(QKV_weight_out_7_14), .input_weight_15(QKV_weight_out_7_15),
                          .input_data_0(QKV_data_out_7_0), .input_data_1(QKV_data_out_7_1), .input_data_2(QKV_data_out_7_2), .input_data_3(QKV_data_out_7_3), .input_data_4(QKV_data_out_7_4), .input_data_5(QKV_data_out_7_5), .input_data_6(QKV_data_out_7_6), .input_data_7(QKV_data_out_7_7), .input_data_8(QKV_data_out_7_8), .input_data_9(QKV_data_out_7_9), .input_data_10(QKV_data_out_7_10), .input_data_11(QKV_data_out_7_11), .input_data_12(QKV_data_out_7_12), .input_data_13(QKV_data_out_7_13), .input_data_14(QKV_data_out_7_14), .input_data_15(QKV_data_out_7_15),
                          .is_write_(QKV_is_write_out_7), .select_(QKV_selcet_out_7),
                          .calc_result_0(QKV_calc_result_7_0), .calc_result_1(QKV_calc_result_7_1), .calc_result_2(QKV_calc_result_7_2), .calc_result_3(QKV_calc_result_7_3), .calc_result_4(QKV_calc_result_7_4), .calc_result_5(QKV_calc_result_7_5), .calc_result_6(QKV_calc_result_7_6), .calc_result_7(QKV_calc_result_7_7), .calc_result_8(QKV_calc_result_7_8), .calc_result_9(QKV_calc_result_7_9), .calc_result_10(QKV_calc_result_7_10), .calc_result_11(QKV_calc_result_7_11), .calc_result_12(QKV_calc_result_7_12), .calc_result_13(QKV_calc_result_7_13), .calc_result_14(QKV_calc_result_7_14), .calc_result_15(QKV_calc_result_7_15)
);

dimc_macro i_dimc_macro_8(.input_addr(QKV_addr_out_8),
                          .input_weight_0(QKV_weight_out_8_0), .input_weight_1(QKV_weight_out_8_1), .input_weight_2(QKV_weight_out_8_2), .input_weight_3(QKV_weight_out_8_3), .input_weight_4(QKV_weight_out_8_4), .input_weight_5(QKV_weight_out_8_5), .input_weight_6(QKV_weight_out_8_6), .input_weight_7(QKV_weight_out_8_7), .input_weight_8(QKV_weight_out_8_8), .input_weight_9(QKV_weight_out_8_9), .input_weight_10(QKV_weight_out_8_10), .input_weight_11(QKV_weight_out_8_11), .input_weight_12(QKV_weight_out_8_12), .input_weight_13(QKV_weight_out_8_13), .input_weight_14(QKV_weight_out_8_14), .input_weight_15(QKV_weight_out_8_15),
                          .input_data_0(QKV_data_out_8_0), .input_data_1(QKV_data_out_8_1), .input_data_2(QKV_data_out_8_2), .input_data_3(QKV_data_out_8_3), .input_data_4(QKV_data_out_8_4), .input_data_5(QKV_data_out_8_5), .input_data_6(QKV_data_out_8_6), .input_data_7(QKV_data_out_8_7), .input_data_8(QKV_data_out_8_8), .input_data_9(QKV_data_out_8_9), .input_data_10(QKV_data_out_8_10), .input_data_11(QKV_data_out_8_11), .input_data_12(QKV_data_out_8_12), .input_data_13(QKV_data_out_8_13), .input_data_14(QKV_data_out_8_14), .input_data_15(QKV_data_out_8_15),
                          .is_write_(QKV_is_write_out_8), .select_(QKV_selcet_out_8),
                          .calc_result_0(QKV_calc_result_8_0), .calc_result_1(QKV_calc_result_8_1), .calc_result_2(QKV_calc_result_8_2), .calc_result_3(QKV_calc_result_8_3), .calc_result_4(QKV_calc_result_8_4), .calc_result_5(QKV_calc_result_8_5), .calc_result_6(QKV_calc_result_8_6), .calc_result_7(QKV_calc_result_8_7), .calc_result_8(QKV_calc_result_8_8), .calc_result_9(QKV_calc_result_8_9), .calc_result_10(QKV_calc_result_8_10), .calc_result_11(QKV_calc_result_8_11), .calc_result_12(QKV_calc_result_8_12), .calc_result_13(QKV_calc_result_8_13), .calc_result_14(QKV_calc_result_8_14), .calc_result_15(QKV_calc_result_8_15)
);

dimc_macro i_dimc_macro_9(.input_addr(QKV_addr_out_9),
                          .input_weight_0(QKV_weight_out_9_0), .input_weight_1(QKV_weight_out_9_1), .input_weight_2(QKV_weight_out_9_2), .input_weight_3(QKV_weight_out_9_3), .input_weight_4(QKV_weight_out_9_4), .input_weight_5(QKV_weight_out_9_5), .input_weight_6(QKV_weight_out_9_6), .input_weight_7(QKV_weight_out_9_7), .input_weight_8(QKV_weight_out_9_8), .input_weight_9(QKV_weight_out_9_9), .input_weight_10(QKV_weight_out_9_10), .input_weight_11(QKV_weight_out_9_11), .input_weight_12(QKV_weight_out_9_12), .input_weight_13(QKV_weight_out_9_13), .input_weight_14(QKV_weight_out_9_14), .input_weight_15(QKV_weight_out_9_15),
                          .input_data_0(QKV_data_out_9_0), .input_data_1(QKV_data_out_9_1), .input_data_2(QKV_data_out_9_2), .input_data_3(QKV_data_out_9_3), .input_data_4(QKV_data_out_9_4), .input_data_5(QKV_data_out_9_5), .input_data_6(QKV_data_out_9_6), .input_data_7(QKV_data_out_9_7), .input_data_8(QKV_data_out_9_8), .input_data_9(QKV_data_out_9_9), .input_data_10(QKV_data_out_9_10), .input_data_11(QKV_data_out_9_11), .input_data_12(QKV_data_out_9_12), .input_data_13(QKV_data_out_9_13), .input_data_14(QKV_data_out_9_14), .input_data_15(QKV_data_out_9_15),
                          .is_write_(QKV_is_write_out_9), .select_(QKV_selcet_out_9),
                          .calc_result_0(QKV_calc_result_9_0), .calc_result_1(QKV_calc_result_9_1), .calc_result_2(QKV_calc_result_9_2), .calc_result_3(QKV_calc_result_9_3), .calc_result_4(QKV_calc_result_9_4), .calc_result_5(QKV_calc_result_9_5), .calc_result_6(QKV_calc_result_9_6), .calc_result_7(QKV_calc_result_9_7), .calc_result_8(QKV_calc_result_9_8), .calc_result_9(QKV_calc_result_9_9), .calc_result_10(QKV_calc_result_9_10), .calc_result_11(QKV_calc_result_9_11), .calc_result_12(QKV_calc_result_9_12), .calc_result_13(QKV_calc_result_9_13), .calc_result_14(QKV_calc_result_9_14), .calc_result_15(QKV_calc_result_9_15)
);

dimc_macro i_dimc_macro_10(.input_addr(QKV_addr_out_10),
                          .input_weight_0(QKV_weight_out_10_0), .input_weight_1(QKV_weight_out_10_1), .input_weight_2(QKV_weight_out_10_2), .input_weight_3(QKV_weight_out_10_3), .input_weight_4(QKV_weight_out_10_4), .input_weight_5(QKV_weight_out_10_5), .input_weight_6(QKV_weight_out_10_6), .input_weight_7(QKV_weight_out_10_7), .input_weight_8(QKV_weight_out_10_8), .input_weight_9(QKV_weight_out_10_9), .input_weight_10(QKV_weight_out_10_10), .input_weight_11(QKV_weight_out_10_11), .input_weight_12(QKV_weight_out_10_12), .input_weight_13(QKV_weight_out_10_13), .input_weight_14(QKV_weight_out_10_14), .input_weight_15(QKV_weight_out_10_15),
                          .input_data_0(QKV_data_out_10_0), .input_data_1(QKV_data_out_10_1), .input_data_2(QKV_data_out_10_2), .input_data_3(QKV_data_out_10_3), .input_data_4(QKV_data_out_10_4), .input_data_5(QKV_data_out_10_5), .input_data_6(QKV_data_out_10_6), .input_data_7(QKV_data_out_10_7), .input_data_8(QKV_data_out_10_8), .input_data_9(QKV_data_out_10_9), .input_data_10(QKV_data_out_10_10), .input_data_11(QKV_data_out_10_11), .input_data_12(QKV_data_out_10_12), .input_data_13(QKV_data_out_10_13), .input_data_14(QKV_data_out_10_14), .input_data_15(QKV_data_out_10_15),
                          .is_write_(QKV_is_write_out_10), .select_(QKV_selcet_out_10),
                          .calc_result_0(QKV_calc_result_10_0), .calc_result_1(QKV_calc_result_10_1), .calc_result_2(QKV_calc_result_10_2), .calc_result_3(QKV_calc_result_10_3), .calc_result_4(QKV_calc_result_10_4), .calc_result_5(QKV_calc_result_10_5), .calc_result_6(QKV_calc_result_10_6), .calc_result_7(QKV_calc_result_10_7), .calc_result_8(QKV_calc_result_10_8), .calc_result_9(QKV_calc_result_10_9), .calc_result_10(QKV_calc_result_10_10), .calc_result_11(QKV_calc_result_10_11), .calc_result_12(QKV_calc_result_10_12), .calc_result_13(QKV_calc_result_10_13), .calc_result_14(QKV_calc_result_10_14), .calc_result_15(QKV_calc_result_10_15)
);

dimc_macro i_dimc_macro_11(.input_addr(QKV_addr_out_11),
                          .input_weight_0(QKV_weight_out_11_0), .input_weight_1(QKV_weight_out_11_1), .input_weight_2(QKV_weight_out_11_2), .input_weight_3(QKV_weight_out_11_3), .input_weight_4(QKV_weight_out_11_4), .input_weight_5(QKV_weight_out_11_5), .input_weight_6(QKV_weight_out_11_6), .input_weight_7(QKV_weight_out_11_7), .input_weight_8(QKV_weight_out_11_8), .input_weight_9(QKV_weight_out_11_9), .input_weight_10(QKV_weight_out_11_10), .input_weight_11(QKV_weight_out_11_11), .input_weight_12(QKV_weight_out_11_12), .input_weight_13(QKV_weight_out_11_13), .input_weight_14(QKV_weight_out_11_14), .input_weight_15(QKV_weight_out_11_15),
                          .input_data_0(QKV_data_out_11_0), .input_data_1(QKV_data_out_11_1), .input_data_2(QKV_data_out_11_2), .input_data_3(QKV_data_out_11_3), .input_data_4(QKV_data_out_11_4), .input_data_5(QKV_data_out_11_5), .input_data_6(QKV_data_out_11_6), .input_data_7(QKV_data_out_11_7), .input_data_8(QKV_data_out_11_8), .input_data_9(QKV_data_out_11_9), .input_data_10(QKV_data_out_11_10), .input_data_11(QKV_data_out_11_11), .input_data_12(QKV_data_out_11_12), .input_data_13(QKV_data_out_11_13), .input_data_14(QKV_data_out_11_14), .input_data_15(QKV_data_out_11_15),
                          .is_write_(QKV_is_write_out_11), .select_(QKV_selcet_out_11),
                          .calc_result_0(QKV_calc_result_11_0), .calc_result_1(QKV_calc_result_11_1), .calc_result_2(QKV_calc_result_11_2), .calc_result_3(QKV_calc_result_11_3), .calc_result_4(QKV_calc_result_11_4), .calc_result_5(QKV_calc_result_11_5), .calc_result_6(QKV_calc_result_11_6), .calc_result_7(QKV_calc_result_11_7), .calc_result_8(QKV_calc_result_11_8), .calc_result_9(QKV_calc_result_11_9), .calc_result_10(QKV_calc_result_11_10), .calc_result_11(QKV_calc_result_11_11), .calc_result_12(QKV_calc_result_11_12), .calc_result_13(QKV_calc_result_11_13), .calc_result_14(QKV_calc_result_11_14), .calc_result_15(QKV_calc_result_11_15)
);

dimc_macro i_dimc_macro_12(.input_addr(QKV_addr_out_12),
                          .input_weight_0(QKV_weight_out_12_0), .input_weight_1(QKV_weight_out_12_1), .input_weight_2(QKV_weight_out_12_2), .input_weight_3(QKV_weight_out_12_3), .input_weight_4(QKV_weight_out_12_4), .input_weight_5(QKV_weight_out_12_5), .input_weight_6(QKV_weight_out_12_6), .input_weight_7(QKV_weight_out_12_7), .input_weight_8(QKV_weight_out_12_8), .input_weight_9(QKV_weight_out_12_9), .input_weight_10(QKV_weight_out_12_10), .input_weight_11(QKV_weight_out_12_11), .input_weight_12(QKV_weight_out_12_12), .input_weight_13(QKV_weight_out_12_13), .input_weight_14(QKV_weight_out_12_14), .input_weight_15(QKV_weight_out_12_15),
                          .input_data_0(QKV_data_out_12_0), .input_data_1(QKV_data_out_12_1), .input_data_2(QKV_data_out_12_2), .input_data_3(QKV_data_out_12_3), .input_data_4(QKV_data_out_12_4), .input_data_5(QKV_data_out_12_5), .input_data_6(QKV_data_out_12_6), .input_data_7(QKV_data_out_12_7), .input_data_8(QKV_data_out_12_8), .input_data_9(QKV_data_out_12_9), .input_data_10(QKV_data_out_12_10), .input_data_11(QKV_data_out_12_11), .input_data_12(QKV_data_out_12_12), .input_data_13(QKV_data_out_12_13), .input_data_14(QKV_data_out_12_14), .input_data_15(QKV_data_out_12_15),
                          .is_write_(QKV_is_write_out_12), .select_(QKV_selcet_out_12),
                          .calc_result_0(QKV_calc_result_12_0), .calc_result_1(QKV_calc_result_12_1), .calc_result_2(QKV_calc_result_12_2), .calc_result_3(QKV_calc_result_12_3), .calc_result_4(QKV_calc_result_12_4), .calc_result_5(QKV_calc_result_12_5), .calc_result_6(QKV_calc_result_12_6), .calc_result_7(QKV_calc_result_12_7), .calc_result_8(QKV_calc_result_12_8), .calc_result_9(QKV_calc_result_12_9), .calc_result_10(QKV_calc_result_12_10), .calc_result_11(QKV_calc_result_12_11), .calc_result_12(QKV_calc_result_12_12), .calc_result_13(QKV_calc_result_12_13), .calc_result_14(QKV_calc_result_12_14), .calc_result_15(QKV_calc_result_12_15)
);

dimc_macro i_dimc_macro_13(.input_addr(QKV_addr_out_13),
                          .input_weight_0(QKV_weight_out_13_0), .input_weight_1(QKV_weight_out_13_1), .input_weight_2(QKV_weight_out_13_2), .input_weight_3(QKV_weight_out_13_3), .input_weight_4(QKV_weight_out_13_4), .input_weight_5(QKV_weight_out_13_5), .input_weight_6(QKV_weight_out_13_6), .input_weight_7(QKV_weight_out_13_7), .input_weight_8(QKV_weight_out_13_8), .input_weight_9(QKV_weight_out_13_9), .input_weight_10(QKV_weight_out_13_10), .input_weight_11(QKV_weight_out_13_11), .input_weight_12(QKV_weight_out_13_12), .input_weight_13(QKV_weight_out_13_13), .input_weight_14(QKV_weight_out_13_14), .input_weight_15(QKV_weight_out_13_15),
                          .input_data_0(QKV_data_out_13_0), .input_data_1(QKV_data_out_13_1), .input_data_2(QKV_data_out_13_2), .input_data_3(QKV_data_out_13_3), .input_data_4(QKV_data_out_13_4), .input_data_5(QKV_data_out_13_5), .input_data_6(QKV_data_out_13_6), .input_data_7(QKV_data_out_13_7), .input_data_8(QKV_data_out_13_8), .input_data_9(QKV_data_out_13_9), .input_data_10(QKV_data_out_13_10), .input_data_11(QKV_data_out_13_11), .input_data_12(QKV_data_out_13_12), .input_data_13(QKV_data_out_13_13), .input_data_14(QKV_data_out_13_14), .input_data_15(QKV_data_out_13_15),
                          .is_write_(QKV_is_write_out_13), .select_(QKV_selcet_out_13),
                          .calc_result_0(QKV_calc_result_13_0), .calc_result_1(QKV_calc_result_13_1), .calc_result_2(QKV_calc_result_13_2), .calc_result_3(QKV_calc_result_13_3), .calc_result_4(QKV_calc_result_13_4), .calc_result_5(QKV_calc_result_13_5), .calc_result_6(QKV_calc_result_13_6), .calc_result_7(QKV_calc_result_13_7), .calc_result_8(QKV_calc_result_13_8), .calc_result_9(QKV_calc_result_13_9), .calc_result_10(QKV_calc_result_13_10), .calc_result_11(QKV_calc_result_13_11), .calc_result_12(QKV_calc_result_13_12), .calc_result_13(QKV_calc_result_13_13), .calc_result_14(QKV_calc_result_13_14), .calc_result_15(QKV_calc_result_13_15)
);

dimc_macro i_dimc_macro_14(.input_addr(QKV_addr_out_14),
                          .input_weight_0(QKV_weight_out_14_0), .input_weight_1(QKV_weight_out_14_1), .input_weight_2(QKV_weight_out_14_2), .input_weight_3(QKV_weight_out_14_3), .input_weight_4(QKV_weight_out_14_4), .input_weight_5(QKV_weight_out_14_5), .input_weight_6(QKV_weight_out_14_6), .input_weight_7(QKV_weight_out_14_7), .input_weight_8(QKV_weight_out_14_8), .input_weight_9(QKV_weight_out_14_9), .input_weight_10(QKV_weight_out_14_10), .input_weight_11(QKV_weight_out_14_11), .input_weight_12(QKV_weight_out_14_12), .input_weight_13(QKV_weight_out_14_13), .input_weight_14(QKV_weight_out_14_14), .input_weight_15(QKV_weight_out_14_15),
                          .input_data_0(QKV_data_out_14_0), .input_data_1(QKV_data_out_14_1), .input_data_2(QKV_data_out_14_2), .input_data_3(QKV_data_out_14_3), .input_data_4(QKV_data_out_14_4), .input_data_5(QKV_data_out_14_5), .input_data_6(QKV_data_out_14_6), .input_data_7(QKV_data_out_14_7), .input_data_8(QKV_data_out_14_8), .input_data_9(QKV_data_out_14_9), .input_data_10(QKV_data_out_14_10), .input_data_11(QKV_data_out_14_11), .input_data_12(QKV_data_out_14_12), .input_data_13(QKV_data_out_14_13), .input_data_14(QKV_data_out_14_14), .input_data_15(QKV_data_out_14_15),
                          .is_write_(QKV_is_write_out_14), .select_(QKV_selcet_out_14),
                          .calc_result_0(QKV_calc_result_14_0), .calc_result_1(QKV_calc_result_14_1), .calc_result_2(QKV_calc_result_14_2), .calc_result_3(QKV_calc_result_14_3), .calc_result_4(QKV_calc_result_14_4), .calc_result_5(QKV_calc_result_14_5), .calc_result_6(QKV_calc_result_14_6), .calc_result_7(QKV_calc_result_14_7), .calc_result_8(QKV_calc_result_14_8), .calc_result_9(QKV_calc_result_14_9), .calc_result_10(QKV_calc_result_14_10), .calc_result_11(QKV_calc_result_14_11), .calc_result_12(QKV_calc_result_14_12), .calc_result_13(QKV_calc_result_14_13), .calc_result_14(QKV_calc_result_14_14), .calc_result_15(QKV_calc_result_14_15)
);

dimc_macro i_dimc_macro_15(.input_addr(QKV_addr_out_15),
                          .input_weight_0(QKV_weight_out_15_0), .input_weight_1(QKV_weight_out_15_1), .input_weight_2(QKV_weight_out_15_2), .input_weight_3(QKV_weight_out_15_3), .input_weight_4(QKV_weight_out_15_4), .input_weight_5(QKV_weight_out_15_5), .input_weight_6(QKV_weight_out_15_6), .input_weight_7(QKV_weight_out_15_7), .input_weight_8(QKV_weight_out_15_8), .input_weight_9(QKV_weight_out_15_9), .input_weight_10(QKV_weight_out_15_10), .input_weight_11(QKV_weight_out_15_11), .input_weight_12(QKV_weight_out_15_12), .input_weight_13(QKV_weight_out_15_13), .input_weight_14(QKV_weight_out_15_14), .input_weight_15(QKV_weight_out_15_15),
                          .input_data_0(QKV_data_out_15_0), .input_data_1(QKV_data_out_15_1), .input_data_2(QKV_data_out_15_2), .input_data_3(QKV_data_out_15_3), .input_data_4(QKV_data_out_15_4), .input_data_5(QKV_data_out_15_5), .input_data_6(QKV_data_out_15_6), .input_data_7(QKV_data_out_15_7), .input_data_8(QKV_data_out_15_8), .input_data_9(QKV_data_out_15_9), .input_data_10(QKV_data_out_15_10), .input_data_11(QKV_data_out_15_11), .input_data_12(QKV_data_out_15_12), .input_data_13(QKV_data_out_15_13), .input_data_14(QKV_data_out_15_14), .input_data_15(QKV_data_out_15_15),
                          .is_write_(QKV_is_write_out_15), .select_(QKV_selcet_out_15),
                          .calc_result_0(QKV_calc_result_15_0), .calc_result_1(QKV_calc_result_15_1), .calc_result_2(QKV_calc_result_15_2), .calc_result_3(QKV_calc_result_15_3), .calc_result_4(QKV_calc_result_15_4), .calc_result_5(QKV_calc_result_15_5), .calc_result_6(QKV_calc_result_15_6), .calc_result_7(QKV_calc_result_15_7), .calc_result_8(QKV_calc_result_15_8), .calc_result_9(QKV_calc_result_15_9), .calc_result_10(QKV_calc_result_15_10), .calc_result_11(QKV_calc_result_15_11), .calc_result_12(QKV_calc_result_15_12), .calc_result_13(QKV_calc_result_15_13), .calc_result_14(QKV_calc_result_15_14), .calc_result_15(QKV_calc_result_15_15)
);

dimc_macro i_dimc_macro_16(.input_addr(QKV_addr_out_16),
                          .input_weight_0(QKV_weight_out_16_0), .input_weight_1(QKV_weight_out_16_1), .input_weight_2(QKV_weight_out_16_2), .input_weight_3(QKV_weight_out_16_3), .input_weight_4(QKV_weight_out_16_4), .input_weight_5(QKV_weight_out_16_5), .input_weight_6(QKV_weight_out_16_6), .input_weight_7(QKV_weight_out_16_7), .input_weight_8(QKV_weight_out_16_8), .input_weight_9(QKV_weight_out_16_9), .input_weight_10(QKV_weight_out_16_10), .input_weight_11(QKV_weight_out_16_11), .input_weight_12(QKV_weight_out_16_12), .input_weight_13(QKV_weight_out_16_13), .input_weight_14(QKV_weight_out_16_14), .input_weight_15(QKV_weight_out_16_15),
                          .input_data_0(QKV_data_out_16_0), .input_data_1(QKV_data_out_16_1), .input_data_2(QKV_data_out_16_2), .input_data_3(QKV_data_out_16_3), .input_data_4(QKV_data_out_16_4), .input_data_5(QKV_data_out_16_5), .input_data_6(QKV_data_out_16_6), .input_data_7(QKV_data_out_16_7), .input_data_8(QKV_data_out_16_8), .input_data_9(QKV_data_out_16_9), .input_data_10(QKV_data_out_16_10), .input_data_11(QKV_data_out_16_11), .input_data_12(QKV_data_out_16_12), .input_data_13(QKV_data_out_16_13), .input_data_14(QKV_data_out_16_14), .input_data_15(QKV_data_out_16_15),
                          .is_write_(QKV_is_write_out_16), .select_(QKV_selcet_out_16),
                          .calc_result_0(QKV_calc_result_16_0), .calc_result_1(QKV_calc_result_16_1), .calc_result_2(QKV_calc_result_16_2), .calc_result_3(QKV_calc_result_16_3), .calc_result_4(QKV_calc_result_16_4), .calc_result_5(QKV_calc_result_16_5), .calc_result_6(QKV_calc_result_16_6), .calc_result_7(QKV_calc_result_16_7), .calc_result_8(QKV_calc_result_16_8), .calc_result_9(QKV_calc_result_16_9), .calc_result_10(QKV_calc_result_16_10), .calc_result_11(QKV_calc_result_16_11), .calc_result_12(QKV_calc_result_16_12), .calc_result_13(QKV_calc_result_16_13), .calc_result_14(QKV_calc_result_16_14), .calc_result_15(QKV_calc_result_16_15)
);

dimc_macro i_dimc_macro_17(.input_addr(QKV_addr_out_17),
                          .input_weight_0(QKV_weight_out_17_0), .input_weight_1(QKV_weight_out_17_1), .input_weight_2(QKV_weight_out_17_2), .input_weight_3(QKV_weight_out_17_3), .input_weight_4(QKV_weight_out_17_4), .input_weight_5(QKV_weight_out_17_5), .input_weight_6(QKV_weight_out_17_6), .input_weight_7(QKV_weight_out_17_7), .input_weight_8(QKV_weight_out_17_8), .input_weight_9(QKV_weight_out_17_9), .input_weight_10(QKV_weight_out_17_10), .input_weight_11(QKV_weight_out_17_11), .input_weight_12(QKV_weight_out_17_12), .input_weight_13(QKV_weight_out_17_13), .input_weight_14(QKV_weight_out_17_14), .input_weight_15(QKV_weight_out_17_15),
                          .input_data_0(QKV_data_out_17_0), .input_data_1(QKV_data_out_17_1), .input_data_2(QKV_data_out_17_2), .input_data_3(QKV_data_out_17_3), .input_data_4(QKV_data_out_17_4), .input_data_5(QKV_data_out_17_5), .input_data_6(QKV_data_out_17_6), .input_data_7(QKV_data_out_17_7), .input_data_8(QKV_data_out_17_8), .input_data_9(QKV_data_out_17_9), .input_data_10(QKV_data_out_17_10), .input_data_11(QKV_data_out_17_11), .input_data_12(QKV_data_out_17_12), .input_data_13(QKV_data_out_17_13), .input_data_14(QKV_data_out_17_14), .input_data_15(QKV_data_out_17_15),
                          .is_write_(QKV_is_write_out_17), .select_(QKV_selcet_out_17),
                          .calc_result_0(QKV_calc_result_17_0), .calc_result_1(QKV_calc_result_17_1), .calc_result_2(QKV_calc_result_17_2), .calc_result_3(QKV_calc_result_17_3), .calc_result_4(QKV_calc_result_17_4), .calc_result_5(QKV_calc_result_17_5), .calc_result_6(QKV_calc_result_17_6), .calc_result_7(QKV_calc_result_17_7), .calc_result_8(QKV_calc_result_17_8), .calc_result_9(QKV_calc_result_17_9), .calc_result_10(QKV_calc_result_17_10), .calc_result_11(QKV_calc_result_17_11), .calc_result_12(QKV_calc_result_17_12), .calc_result_13(QKV_calc_result_17_13), .calc_result_14(QKV_calc_result_17_14), .calc_result_15(QKV_calc_result_17_15)
);

dimc_macro i_dimc_macro_18(.input_addr(QKV_addr_out_18),
                          .input_weight_0(QKV_weight_out_18_0), .input_weight_1(QKV_weight_out_18_1), .input_weight_2(QKV_weight_out_18_2), .input_weight_3(QKV_weight_out_18_3), .input_weight_4(QKV_weight_out_18_4), .input_weight_5(QKV_weight_out_18_5), .input_weight_6(QKV_weight_out_18_6), .input_weight_7(QKV_weight_out_18_7), .input_weight_8(QKV_weight_out_18_8), .input_weight_9(QKV_weight_out_18_9), .input_weight_10(QKV_weight_out_18_10), .input_weight_11(QKV_weight_out_18_11), .input_weight_12(QKV_weight_out_18_12), .input_weight_13(QKV_weight_out_18_13), .input_weight_14(QKV_weight_out_18_14), .input_weight_15(QKV_weight_out_18_15),
                          .input_data_0(QKV_data_out_18_0), .input_data_1(QKV_data_out_18_1), .input_data_2(QKV_data_out_18_2), .input_data_3(QKV_data_out_18_3), .input_data_4(QKV_data_out_18_4), .input_data_5(QKV_data_out_18_5), .input_data_6(QKV_data_out_18_6), .input_data_7(QKV_data_out_18_7), .input_data_8(QKV_data_out_18_8), .input_data_9(QKV_data_out_18_9), .input_data_10(QKV_data_out_18_10), .input_data_11(QKV_data_out_18_11), .input_data_12(QKV_data_out_18_12), .input_data_13(QKV_data_out_18_13), .input_data_14(QKV_data_out_18_14), .input_data_15(QKV_data_out_18_15),
                          .is_write_(QKV_is_write_out_18), .select_(QKV_selcet_out_18),
                          .calc_result_0(QKV_calc_result_18_0), .calc_result_1(QKV_calc_result_18_1), .calc_result_2(QKV_calc_result_18_2), .calc_result_3(QKV_calc_result_18_3), .calc_result_4(QKV_calc_result_18_4), .calc_result_5(QKV_calc_result_18_5), .calc_result_6(QKV_calc_result_18_6), .calc_result_7(QKV_calc_result_18_7), .calc_result_8(QKV_calc_result_18_8), .calc_result_9(QKV_calc_result_18_9), .calc_result_10(QKV_calc_result_18_10), .calc_result_11(QKV_calc_result_18_11), .calc_result_12(QKV_calc_result_18_12), .calc_result_13(QKV_calc_result_18_13), .calc_result_14(QKV_calc_result_18_14), .calc_result_15(QKV_calc_result_18_15)
);

dimc_macro i_dimc_macro_19(.input_addr(QKV_addr_out_19),
                          .input_weight_0(QKV_weight_out_19_0), .input_weight_1(QKV_weight_out_19_1), .input_weight_2(QKV_weight_out_19_2), .input_weight_3(QKV_weight_out_19_3), .input_weight_4(QKV_weight_out_19_4), .input_weight_5(QKV_weight_out_19_5), .input_weight_6(QKV_weight_out_19_6), .input_weight_7(QKV_weight_out_19_7), .input_weight_8(QKV_weight_out_19_8), .input_weight_9(QKV_weight_out_19_9), .input_weight_10(QKV_weight_out_19_10), .input_weight_11(QKV_weight_out_19_11), .input_weight_12(QKV_weight_out_19_12), .input_weight_13(QKV_weight_out_19_13), .input_weight_14(QKV_weight_out_19_14), .input_weight_15(QKV_weight_out_19_15),
                          .input_data_0(QKV_data_out_19_0), .input_data_1(QKV_data_out_19_1), .input_data_2(QKV_data_out_19_2), .input_data_3(QKV_data_out_19_3), .input_data_4(QKV_data_out_19_4), .input_data_5(QKV_data_out_19_5), .input_data_6(QKV_data_out_19_6), .input_data_7(QKV_data_out_19_7), .input_data_8(QKV_data_out_19_8), .input_data_9(QKV_data_out_19_9), .input_data_10(QKV_data_out_19_10), .input_data_11(QKV_data_out_19_11), .input_data_12(QKV_data_out_19_12), .input_data_13(QKV_data_out_19_13), .input_data_14(QKV_data_out_19_14), .input_data_15(QKV_data_out_19_15),
                          .is_write_(QKV_is_write_out_19), .select_(QKV_selcet_out_19),
                          .calc_result_0(QKV_calc_result_19_0), .calc_result_1(QKV_calc_result_19_1), .calc_result_2(QKV_calc_result_19_2), .calc_result_3(QKV_calc_result_19_3), .calc_result_4(QKV_calc_result_19_4), .calc_result_5(QKV_calc_result_19_5), .calc_result_6(QKV_calc_result_19_6), .calc_result_7(QKV_calc_result_19_7), .calc_result_8(QKV_calc_result_19_8), .calc_result_9(QKV_calc_result_19_9), .calc_result_10(QKV_calc_result_19_10), .calc_result_11(QKV_calc_result_19_11), .calc_result_12(QKV_calc_result_19_12), .calc_result_13(QKV_calc_result_19_13), .calc_result_14(QKV_calc_result_19_14), .calc_result_15(QKV_calc_result_19_15)
);

dimc_macro i_dimc_macro_20(.input_addr(QKV_addr_out_20),
                          .input_weight_0(QKV_weight_out_20_0), .input_weight_1(QKV_weight_out_20_1), .input_weight_2(QKV_weight_out_20_2), .input_weight_3(QKV_weight_out_20_3), .input_weight_4(QKV_weight_out_20_4), .input_weight_5(QKV_weight_out_20_5), .input_weight_6(QKV_weight_out_20_6), .input_weight_7(QKV_weight_out_20_7), .input_weight_8(QKV_weight_out_20_8), .input_weight_9(QKV_weight_out_20_9), .input_weight_10(QKV_weight_out_20_10), .input_weight_11(QKV_weight_out_20_11), .input_weight_12(QKV_weight_out_20_12), .input_weight_13(QKV_weight_out_20_13), .input_weight_14(QKV_weight_out_20_14), .input_weight_15(QKV_weight_out_20_15),
                          .input_data_0(QKV_data_out_20_0), .input_data_1(QKV_data_out_20_1), .input_data_2(QKV_data_out_20_2), .input_data_3(QKV_data_out_20_3), .input_data_4(QKV_data_out_20_4), .input_data_5(QKV_data_out_20_5), .input_data_6(QKV_data_out_20_6), .input_data_7(QKV_data_out_20_7), .input_data_8(QKV_data_out_20_8), .input_data_9(QKV_data_out_20_9), .input_data_10(QKV_data_out_20_10), .input_data_11(QKV_data_out_20_11), .input_data_12(QKV_data_out_20_12), .input_data_13(QKV_data_out_20_13), .input_data_14(QKV_data_out_20_14), .input_data_15(QKV_data_out_20_15),
                          .is_write_(QKV_is_write_out_20), .select_(QKV_selcet_out_20),
                          .calc_result_0(QKV_calc_result_20_0), .calc_result_1(QKV_calc_result_20_1), .calc_result_2(QKV_calc_result_20_2), .calc_result_3(QKV_calc_result_20_3), .calc_result_4(QKV_calc_result_20_4), .calc_result_5(QKV_calc_result_20_5), .calc_result_6(QKV_calc_result_20_6), .calc_result_7(QKV_calc_result_20_7), .calc_result_8(QKV_calc_result_20_8), .calc_result_9(QKV_calc_result_20_9), .calc_result_10(QKV_calc_result_20_10), .calc_result_11(QKV_calc_result_20_11), .calc_result_12(QKV_calc_result_20_12), .calc_result_13(QKV_calc_result_20_13), .calc_result_14(QKV_calc_result_20_14), .calc_result_15(QKV_calc_result_20_15)
);

dimc_macro i_dimc_macro_21(.input_addr(QKV_addr_out_21),
                          .input_weight_0(QKV_weight_out_21_0), .input_weight_1(QKV_weight_out_21_1), .input_weight_2(QKV_weight_out_21_2), .input_weight_3(QKV_weight_out_21_3), .input_weight_4(QKV_weight_out_21_4), .input_weight_5(QKV_weight_out_21_5), .input_weight_6(QKV_weight_out_21_6), .input_weight_7(QKV_weight_out_21_7), .input_weight_8(QKV_weight_out_21_8), .input_weight_9(QKV_weight_out_21_9), .input_weight_10(QKV_weight_out_21_10), .input_weight_11(QKV_weight_out_21_11), .input_weight_12(QKV_weight_out_21_12), .input_weight_13(QKV_weight_out_21_13), .input_weight_14(QKV_weight_out_21_14), .input_weight_15(QKV_weight_out_21_15),
                          .input_data_0(QKV_data_out_21_0), .input_data_1(QKV_data_out_21_1), .input_data_2(QKV_data_out_21_2), .input_data_3(QKV_data_out_21_3), .input_data_4(QKV_data_out_21_4), .input_data_5(QKV_data_out_21_5), .input_data_6(QKV_data_out_21_6), .input_data_7(QKV_data_out_21_7), .input_data_8(QKV_data_out_21_8), .input_data_9(QKV_data_out_21_9), .input_data_10(QKV_data_out_21_10), .input_data_11(QKV_data_out_21_11), .input_data_12(QKV_data_out_21_12), .input_data_13(QKV_data_out_21_13), .input_data_14(QKV_data_out_21_14), .input_data_15(QKV_data_out_21_15),
                          .is_write_(QKV_is_write_out_21), .select_(QKV_selcet_out_21),
                          .calc_result_0(QKV_calc_result_21_0), .calc_result_1(QKV_calc_result_21_1), .calc_result_2(QKV_calc_result_21_2), .calc_result_3(QKV_calc_result_21_3), .calc_result_4(QKV_calc_result_21_4), .calc_result_5(QKV_calc_result_21_5), .calc_result_6(QKV_calc_result_21_6), .calc_result_7(QKV_calc_result_21_7), .calc_result_8(QKV_calc_result_21_8), .calc_result_9(QKV_calc_result_21_9), .calc_result_10(QKV_calc_result_21_10), .calc_result_11(QKV_calc_result_21_11), .calc_result_12(QKV_calc_result_21_12), .calc_result_13(QKV_calc_result_21_13), .calc_result_14(QKV_calc_result_21_14), .calc_result_15(QKV_calc_result_21_15)
);

dimc_macro i_dimc_macro_22(.input_addr(QKV_addr_out_22),
                          .input_weight_0(QKV_weight_out_22_0), .input_weight_1(QKV_weight_out_22_1), .input_weight_2(QKV_weight_out_22_2), .input_weight_3(QKV_weight_out_22_3), .input_weight_4(QKV_weight_out_22_4), .input_weight_5(QKV_weight_out_22_5), .input_weight_6(QKV_weight_out_22_6), .input_weight_7(QKV_weight_out_22_7), .input_weight_8(QKV_weight_out_22_8), .input_weight_9(QKV_weight_out_22_9), .input_weight_10(QKV_weight_out_22_10), .input_weight_11(QKV_weight_out_22_11), .input_weight_12(QKV_weight_out_22_12), .input_weight_13(QKV_weight_out_22_13), .input_weight_14(QKV_weight_out_22_14), .input_weight_15(QKV_weight_out_22_15),
                          .input_data_0(QKV_data_out_22_0), .input_data_1(QKV_data_out_22_1), .input_data_2(QKV_data_out_22_2), .input_data_3(QKV_data_out_22_3), .input_data_4(QKV_data_out_22_4), .input_data_5(QKV_data_out_22_5), .input_data_6(QKV_data_out_22_6), .input_data_7(QKV_data_out_22_7), .input_data_8(QKV_data_out_22_8), .input_data_9(QKV_data_out_22_9), .input_data_10(QKV_data_out_22_10), .input_data_11(QKV_data_out_22_11), .input_data_12(QKV_data_out_22_12), .input_data_13(QKV_data_out_22_13), .input_data_14(QKV_data_out_22_14), .input_data_15(QKV_data_out_22_15),
                          .is_write_(QKV_is_write_out_22), .select_(QKV_selcet_out_22),
                          .calc_result_0(QKV_calc_result_22_0), .calc_result_1(QKV_calc_result_22_1), .calc_result_2(QKV_calc_result_22_2), .calc_result_3(QKV_calc_result_22_3), .calc_result_4(QKV_calc_result_22_4), .calc_result_5(QKV_calc_result_22_5), .calc_result_6(QKV_calc_result_22_6), .calc_result_7(QKV_calc_result_22_7), .calc_result_8(QKV_calc_result_22_8), .calc_result_9(QKV_calc_result_22_9), .calc_result_10(QKV_calc_result_22_10), .calc_result_11(QKV_calc_result_22_11), .calc_result_12(QKV_calc_result_22_12), .calc_result_13(QKV_calc_result_22_13), .calc_result_14(QKV_calc_result_22_14), .calc_result_15(QKV_calc_result_22_15)
);

dimc_macro i_dimc_macro_23(.input_addr(QKV_addr_out_23),
                          .input_weight_0(QKV_weight_out_23_0), .input_weight_1(QKV_weight_out_23_1), .input_weight_2(QKV_weight_out_23_2), .input_weight_3(QKV_weight_out_23_3), .input_weight_4(QKV_weight_out_23_4), .input_weight_5(QKV_weight_out_23_5), .input_weight_6(QKV_weight_out_23_6), .input_weight_7(QKV_weight_out_23_7), .input_weight_8(QKV_weight_out_23_8), .input_weight_9(QKV_weight_out_23_9), .input_weight_10(QKV_weight_out_23_10), .input_weight_11(QKV_weight_out_23_11), .input_weight_12(QKV_weight_out_23_12), .input_weight_13(QKV_weight_out_23_13), .input_weight_14(QKV_weight_out_23_14), .input_weight_15(QKV_weight_out_23_15),
                          .input_data_0(QKV_data_out_23_0), .input_data_1(QKV_data_out_23_1), .input_data_2(QKV_data_out_23_2), .input_data_3(QKV_data_out_23_3), .input_data_4(QKV_data_out_23_4), .input_data_5(QKV_data_out_23_5), .input_data_6(QKV_data_out_23_6), .input_data_7(QKV_data_out_23_7), .input_data_8(QKV_data_out_23_8), .input_data_9(QKV_data_out_23_9), .input_data_10(QKV_data_out_23_10), .input_data_11(QKV_data_out_23_11), .input_data_12(QKV_data_out_23_12), .input_data_13(QKV_data_out_23_13), .input_data_14(QKV_data_out_23_14), .input_data_15(QKV_data_out_23_15),
                          .is_write_(QKV_is_write_out_23), .select_(QKV_selcet_out_23),
                          .calc_result_0(QKV_calc_result_23_0), .calc_result_1(QKV_calc_result_23_1), .calc_result_2(QKV_calc_result_23_2), .calc_result_3(QKV_calc_result_23_3), .calc_result_4(QKV_calc_result_23_4), .calc_result_5(QKV_calc_result_23_5), .calc_result_6(QKV_calc_result_23_6), .calc_result_7(QKV_calc_result_23_7), .calc_result_8(QKV_calc_result_23_8), .calc_result_9(QKV_calc_result_23_9), .calc_result_10(QKV_calc_result_23_10), .calc_result_11(QKV_calc_result_23_11), .calc_result_12(QKV_calc_result_23_12), .calc_result_13(QKV_calc_result_23_13), .calc_result_14(QKV_calc_result_23_14), .calc_result_15(QKV_calc_result_23_15)
);

dimc_macro i_dimc_macro_24(.input_addr(QKV_addr_out_24),
                          .input_weight_0(QKV_weight_out_24_0), .input_weight_1(QKV_weight_out_24_1), .input_weight_2(QKV_weight_out_24_2), .input_weight_3(QKV_weight_out_24_3), .input_weight_4(QKV_weight_out_24_4), .input_weight_5(QKV_weight_out_24_5), .input_weight_6(QKV_weight_out_24_6), .input_weight_7(QKV_weight_out_24_7), .input_weight_8(QKV_weight_out_24_8), .input_weight_9(QKV_weight_out_24_9), .input_weight_10(QKV_weight_out_24_10), .input_weight_11(QKV_weight_out_24_11), .input_weight_12(QKV_weight_out_24_12), .input_weight_13(QKV_weight_out_24_13), .input_weight_14(QKV_weight_out_24_14), .input_weight_15(QKV_weight_out_24_15),
                          .input_data_0(QKV_data_out_24_0), .input_data_1(QKV_data_out_24_1), .input_data_2(QKV_data_out_24_2), .input_data_3(QKV_data_out_24_3), .input_data_4(QKV_data_out_24_4), .input_data_5(QKV_data_out_24_5), .input_data_6(QKV_data_out_24_6), .input_data_7(QKV_data_out_24_7), .input_data_8(QKV_data_out_24_8), .input_data_9(QKV_data_out_24_9), .input_data_10(QKV_data_out_24_10), .input_data_11(QKV_data_out_24_11), .input_data_12(QKV_data_out_24_12), .input_data_13(QKV_data_out_24_13), .input_data_14(QKV_data_out_24_14), .input_data_15(QKV_data_out_24_15),
                          .is_write_(QKV_is_write_out_24), .select_(QKV_selcet_out_24),
                          .calc_result_0(QKV_calc_result_24_0), .calc_result_1(QKV_calc_result_24_1), .calc_result_2(QKV_calc_result_24_2), .calc_result_3(QKV_calc_result_24_3), .calc_result_4(QKV_calc_result_24_4), .calc_result_5(QKV_calc_result_24_5), .calc_result_6(QKV_calc_result_24_6), .calc_result_7(QKV_calc_result_24_7), .calc_result_8(QKV_calc_result_24_8), .calc_result_9(QKV_calc_result_24_9), .calc_result_10(QKV_calc_result_24_10), .calc_result_11(QKV_calc_result_24_11), .calc_result_12(QKV_calc_result_24_12), .calc_result_13(QKV_calc_result_24_13), .calc_result_14(QKV_calc_result_24_14), .calc_result_15(QKV_calc_result_24_15)
);

dimc_macro i_dimc_macro_25(.input_addr(QKV_addr_out_25),
                          .input_weight_0(QKV_weight_out_25_0), .input_weight_1(QKV_weight_out_25_1), .input_weight_2(QKV_weight_out_25_2), .input_weight_3(QKV_weight_out_25_3), .input_weight_4(QKV_weight_out_25_4), .input_weight_5(QKV_weight_out_25_5), .input_weight_6(QKV_weight_out_25_6), .input_weight_7(QKV_weight_out_25_7), .input_weight_8(QKV_weight_out_25_8), .input_weight_9(QKV_weight_out_25_9), .input_weight_10(QKV_weight_out_25_10), .input_weight_11(QKV_weight_out_25_11), .input_weight_12(QKV_weight_out_25_12), .input_weight_13(QKV_weight_out_25_13), .input_weight_14(QKV_weight_out_25_14), .input_weight_15(QKV_weight_out_25_15),
                          .input_data_0(QKV_data_out_25_0), .input_data_1(QKV_data_out_25_1), .input_data_2(QKV_data_out_25_2), .input_data_3(QKV_data_out_25_3), .input_data_4(QKV_data_out_25_4), .input_data_5(QKV_data_out_25_5), .input_data_6(QKV_data_out_25_6), .input_data_7(QKV_data_out_25_7), .input_data_8(QKV_data_out_25_8), .input_data_9(QKV_data_out_25_9), .input_data_10(QKV_data_out_25_10), .input_data_11(QKV_data_out_25_11), .input_data_12(QKV_data_out_25_12), .input_data_13(QKV_data_out_25_13), .input_data_14(QKV_data_out_25_14), .input_data_15(QKV_data_out_25_15),
                          .is_write_(QKV_is_write_out_25), .select_(QKV_selcet_out_25),
                          .calc_result_0(QKV_calc_result_25_0), .calc_result_1(QKV_calc_result_25_1), .calc_result_2(QKV_calc_result_25_2), .calc_result_3(QKV_calc_result_25_3), .calc_result_4(QKV_calc_result_25_4), .calc_result_5(QKV_calc_result_25_5), .calc_result_6(QKV_calc_result_25_6), .calc_result_7(QKV_calc_result_25_7), .calc_result_8(QKV_calc_result_25_8), .calc_result_9(QKV_calc_result_25_9), .calc_result_10(QKV_calc_result_25_10), .calc_result_11(QKV_calc_result_25_11), .calc_result_12(QKV_calc_result_25_12), .calc_result_13(QKV_calc_result_25_13), .calc_result_14(QKV_calc_result_25_14), .calc_result_15(QKV_calc_result_25_15)
);

dimc_macro i_dimc_macro_26(.input_addr(QKV_addr_out_26),
                          .input_weight_0(QKV_weight_out_26_0), .input_weight_1(QKV_weight_out_26_1), .input_weight_2(QKV_weight_out_26_2), .input_weight_3(QKV_weight_out_26_3), .input_weight_4(QKV_weight_out_26_4), .input_weight_5(QKV_weight_out_26_5), .input_weight_6(QKV_weight_out_26_6), .input_weight_7(QKV_weight_out_26_7), .input_weight_8(QKV_weight_out_26_8), .input_weight_9(QKV_weight_out_26_9), .input_weight_10(QKV_weight_out_26_10), .input_weight_11(QKV_weight_out_26_11), .input_weight_12(QKV_weight_out_26_12), .input_weight_13(QKV_weight_out_26_13), .input_weight_14(QKV_weight_out_26_14), .input_weight_15(QKV_weight_out_26_15),
                          .input_data_0(QKV_data_out_26_0), .input_data_1(QKV_data_out_26_1), .input_data_2(QKV_data_out_26_2), .input_data_3(QKV_data_out_26_3), .input_data_4(QKV_data_out_26_4), .input_data_5(QKV_data_out_26_5), .input_data_6(QKV_data_out_26_6), .input_data_7(QKV_data_out_26_7), .input_data_8(QKV_data_out_26_8), .input_data_9(QKV_data_out_26_9), .input_data_10(QKV_data_out_26_10), .input_data_11(QKV_data_out_26_11), .input_data_12(QKV_data_out_26_12), .input_data_13(QKV_data_out_26_13), .input_data_14(QKV_data_out_26_14), .input_data_15(QKV_data_out_26_15),
                          .is_write_(QKV_is_write_out_26), .select_(QKV_selcet_out_26),
                          .calc_result_0(QKV_calc_result_26_0), .calc_result_1(QKV_calc_result_26_1), .calc_result_2(QKV_calc_result_26_2), .calc_result_3(QKV_calc_result_26_3), .calc_result_4(QKV_calc_result_26_4), .calc_result_5(QKV_calc_result_26_5), .calc_result_6(QKV_calc_result_26_6), .calc_result_7(QKV_calc_result_26_7), .calc_result_8(QKV_calc_result_26_8), .calc_result_9(QKV_calc_result_26_9), .calc_result_10(QKV_calc_result_26_10), .calc_result_11(QKV_calc_result_26_11), .calc_result_12(QKV_calc_result_26_12), .calc_result_13(QKV_calc_result_26_13), .calc_result_14(QKV_calc_result_26_14), .calc_result_15(QKV_calc_result_26_15)
);

dimc_macro i_dimc_macro_27(.input_addr(QKV_addr_out_27),
                          .input_weight_0(QKV_weight_out_27_0), .input_weight_1(QKV_weight_out_27_1), .input_weight_2(QKV_weight_out_27_2), .input_weight_3(QKV_weight_out_27_3), .input_weight_4(QKV_weight_out_27_4), .input_weight_5(QKV_weight_out_27_5), .input_weight_6(QKV_weight_out_27_6), .input_weight_7(QKV_weight_out_27_7), .input_weight_8(QKV_weight_out_27_8), .input_weight_9(QKV_weight_out_27_9), .input_weight_10(QKV_weight_out_27_10), .input_weight_11(QKV_weight_out_27_11), .input_weight_12(QKV_weight_out_27_12), .input_weight_13(QKV_weight_out_27_13), .input_weight_14(QKV_weight_out_27_14), .input_weight_15(QKV_weight_out_27_15),
                          .input_data_0(QKV_data_out_27_0), .input_data_1(QKV_data_out_27_1), .input_data_2(QKV_data_out_27_2), .input_data_3(QKV_data_out_27_3), .input_data_4(QKV_data_out_27_4), .input_data_5(QKV_data_out_27_5), .input_data_6(QKV_data_out_27_6), .input_data_7(QKV_data_out_27_7), .input_data_8(QKV_data_out_27_8), .input_data_9(QKV_data_out_27_9), .input_data_10(QKV_data_out_27_10), .input_data_11(QKV_data_out_27_11), .input_data_12(QKV_data_out_27_12), .input_data_13(QKV_data_out_27_13), .input_data_14(QKV_data_out_27_14), .input_data_15(QKV_data_out_27_15),
                          .is_write_(QKV_is_write_out_27), .select_(QKV_selcet_out_27),
                          .calc_result_0(QKV_calc_result_27_0), .calc_result_1(QKV_calc_result_27_1), .calc_result_2(QKV_calc_result_27_2), .calc_result_3(QKV_calc_result_27_3), .calc_result_4(QKV_calc_result_27_4), .calc_result_5(QKV_calc_result_27_5), .calc_result_6(QKV_calc_result_27_6), .calc_result_7(QKV_calc_result_27_7), .calc_result_8(QKV_calc_result_27_8), .calc_result_9(QKV_calc_result_27_9), .calc_result_10(QKV_calc_result_27_10), .calc_result_11(QKV_calc_result_27_11), .calc_result_12(QKV_calc_result_27_12), .calc_result_13(QKV_calc_result_27_13), .calc_result_14(QKV_calc_result_27_14), .calc_result_15(QKV_calc_result_27_15)
);

dimc_macro i_dimc_macro_28(.input_addr(QKV_addr_out_28),
                          .input_weight_0(QKV_weight_out_28_0), .input_weight_1(QKV_weight_out_28_1), .input_weight_2(QKV_weight_out_28_2), .input_weight_3(QKV_weight_out_28_3), .input_weight_4(QKV_weight_out_28_4), .input_weight_5(QKV_weight_out_28_5), .input_weight_6(QKV_weight_out_28_6), .input_weight_7(QKV_weight_out_28_7), .input_weight_8(QKV_weight_out_28_8), .input_weight_9(QKV_weight_out_28_9), .input_weight_10(QKV_weight_out_28_10), .input_weight_11(QKV_weight_out_28_11), .input_weight_12(QKV_weight_out_28_12), .input_weight_13(QKV_weight_out_28_13), .input_weight_14(QKV_weight_out_28_14), .input_weight_15(QKV_weight_out_28_15),
                          .input_data_0(QKV_data_out_28_0), .input_data_1(QKV_data_out_28_1), .input_data_2(QKV_data_out_28_2), .input_data_3(QKV_data_out_28_3), .input_data_4(QKV_data_out_28_4), .input_data_5(QKV_data_out_28_5), .input_data_6(QKV_data_out_28_6), .input_data_7(QKV_data_out_28_7), .input_data_8(QKV_data_out_28_8), .input_data_9(QKV_data_out_28_9), .input_data_10(QKV_data_out_28_10), .input_data_11(QKV_data_out_28_11), .input_data_12(QKV_data_out_28_12), .input_data_13(QKV_data_out_28_13), .input_data_14(QKV_data_out_28_14), .input_data_15(QKV_data_out_28_15),
                          .is_write_(QKV_is_write_out_28), .select_(QKV_selcet_out_28),
                          .calc_result_0(QKV_calc_result_28_0), .calc_result_1(QKV_calc_result_28_1), .calc_result_2(QKV_calc_result_28_2), .calc_result_3(QKV_calc_result_28_3), .calc_result_4(QKV_calc_result_28_4), .calc_result_5(QKV_calc_result_28_5), .calc_result_6(QKV_calc_result_28_6), .calc_result_7(QKV_calc_result_28_7), .calc_result_8(QKV_calc_result_28_8), .calc_result_9(QKV_calc_result_28_9), .calc_result_10(QKV_calc_result_28_10), .calc_result_11(QKV_calc_result_28_11), .calc_result_12(QKV_calc_result_28_12), .calc_result_13(QKV_calc_result_28_13), .calc_result_14(QKV_calc_result_28_14), .calc_result_15(QKV_calc_result_28_15)
);

dimc_macro i_dimc_macro_29(.input_addr(QKV_addr_out_29),
                          .input_weight_0(QKV_weight_out_29_0), .input_weight_1(QKV_weight_out_29_1), .input_weight_2(QKV_weight_out_29_2), .input_weight_3(QKV_weight_out_29_3), .input_weight_4(QKV_weight_out_29_4), .input_weight_5(QKV_weight_out_29_5), .input_weight_6(QKV_weight_out_29_6), .input_weight_7(QKV_weight_out_29_7), .input_weight_8(QKV_weight_out_29_8), .input_weight_9(QKV_weight_out_29_9), .input_weight_10(QKV_weight_out_29_10), .input_weight_11(QKV_weight_out_29_11), .input_weight_12(QKV_weight_out_29_12), .input_weight_13(QKV_weight_out_29_13), .input_weight_14(QKV_weight_out_29_14), .input_weight_15(QKV_weight_out_29_15),
                          .input_data_0(QKV_data_out_29_0), .input_data_1(QKV_data_out_29_1), .input_data_2(QKV_data_out_29_2), .input_data_3(QKV_data_out_29_3), .input_data_4(QKV_data_out_29_4), .input_data_5(QKV_data_out_29_5), .input_data_6(QKV_data_out_29_6), .input_data_7(QKV_data_out_29_7), .input_data_8(QKV_data_out_29_8), .input_data_9(QKV_data_out_29_9), .input_data_10(QKV_data_out_29_10), .input_data_11(QKV_data_out_29_11), .input_data_12(QKV_data_out_29_12), .input_data_13(QKV_data_out_29_13), .input_data_14(QKV_data_out_29_14), .input_data_15(QKV_data_out_29_15),
                          .is_write_(QKV_is_write_out_29), .select_(QKV_selcet_out_29),
                          .calc_result_0(QKV_calc_result_29_0), .calc_result_1(QKV_calc_result_29_1), .calc_result_2(QKV_calc_result_29_2), .calc_result_3(QKV_calc_result_29_3), .calc_result_4(QKV_calc_result_29_4), .calc_result_5(QKV_calc_result_29_5), .calc_result_6(QKV_calc_result_29_6), .calc_result_7(QKV_calc_result_29_7), .calc_result_8(QKV_calc_result_29_8), .calc_result_9(QKV_calc_result_29_9), .calc_result_10(QKV_calc_result_29_10), .calc_result_11(QKV_calc_result_29_11), .calc_result_12(QKV_calc_result_29_12), .calc_result_13(QKV_calc_result_29_13), .calc_result_14(QKV_calc_result_29_14), .calc_result_15(QKV_calc_result_29_15)
);

dimc_macro i_dimc_macro_30(.input_addr(QKV_addr_out_30),
                          .input_weight_0(QKV_weight_out_30_0), .input_weight_1(QKV_weight_out_30_1), .input_weight_2(QKV_weight_out_30_2), .input_weight_3(QKV_weight_out_30_3), .input_weight_4(QKV_weight_out_30_4), .input_weight_5(QKV_weight_out_30_5), .input_weight_6(QKV_weight_out_30_6), .input_weight_7(QKV_weight_out_30_7), .input_weight_8(QKV_weight_out_30_8), .input_weight_9(QKV_weight_out_30_9), .input_weight_10(QKV_weight_out_30_10), .input_weight_11(QKV_weight_out_30_11), .input_weight_12(QKV_weight_out_30_12), .input_weight_13(QKV_weight_out_30_13), .input_weight_14(QKV_weight_out_30_14), .input_weight_15(QKV_weight_out_30_15),
                          .input_data_0(QKV_data_out_30_0), .input_data_1(QKV_data_out_30_1), .input_data_2(QKV_data_out_30_2), .input_data_3(QKV_data_out_30_3), .input_data_4(QKV_data_out_30_4), .input_data_5(QKV_data_out_30_5), .input_data_6(QKV_data_out_30_6), .input_data_7(QKV_data_out_30_7), .input_data_8(QKV_data_out_30_8), .input_data_9(QKV_data_out_30_9), .input_data_10(QKV_data_out_30_10), .input_data_11(QKV_data_out_30_11), .input_data_12(QKV_data_out_30_12), .input_data_13(QKV_data_out_30_13), .input_data_14(QKV_data_out_30_14), .input_data_15(QKV_data_out_30_15),
                          .is_write_(QKV_is_write_out_30), .select_(QKV_selcet_out_30),
                          .calc_result_0(QKV_calc_result_30_0), .calc_result_1(QKV_calc_result_30_1), .calc_result_2(QKV_calc_result_30_2), .calc_result_3(QKV_calc_result_30_3), .calc_result_4(QKV_calc_result_30_4), .calc_result_5(QKV_calc_result_30_5), .calc_result_6(QKV_calc_result_30_6), .calc_result_7(QKV_calc_result_30_7), .calc_result_8(QKV_calc_result_30_8), .calc_result_9(QKV_calc_result_30_9), .calc_result_10(QKV_calc_result_30_10), .calc_result_11(QKV_calc_result_30_11), .calc_result_12(QKV_calc_result_30_12), .calc_result_13(QKV_calc_result_30_13), .calc_result_14(QKV_calc_result_30_14), .calc_result_15(QKV_calc_result_30_15)
);

dimc_macro i_dimc_macro_31(.input_addr(QKV_addr_out_31),
                          .input_weight_0(QKV_weight_out_31_0), .input_weight_1(QKV_weight_out_31_1), .input_weight_2(QKV_weight_out_31_2), .input_weight_3(QKV_weight_out_31_3), .input_weight_4(QKV_weight_out_31_4), .input_weight_5(QKV_weight_out_31_5), .input_weight_6(QKV_weight_out_31_6), .input_weight_7(QKV_weight_out_31_7), .input_weight_8(QKV_weight_out_31_8), .input_weight_9(QKV_weight_out_31_9), .input_weight_10(QKV_weight_out_31_10), .input_weight_11(QKV_weight_out_31_11), .input_weight_12(QKV_weight_out_31_12), .input_weight_13(QKV_weight_out_31_13), .input_weight_14(QKV_weight_out_31_14), .input_weight_15(QKV_weight_out_31_15),
                          .input_data_0(QKV_data_out_31_0), .input_data_1(QKV_data_out_31_1), .input_data_2(QKV_data_out_31_2), .input_data_3(QKV_data_out_31_3), .input_data_4(QKV_data_out_31_4), .input_data_5(QKV_data_out_31_5), .input_data_6(QKV_data_out_31_6), .input_data_7(QKV_data_out_31_7), .input_data_8(QKV_data_out_31_8), .input_data_9(QKV_data_out_31_9), .input_data_10(QKV_data_out_31_10), .input_data_11(QKV_data_out_31_11), .input_data_12(QKV_data_out_31_12), .input_data_13(QKV_data_out_31_13), .input_data_14(QKV_data_out_31_14), .input_data_15(QKV_data_out_31_15),
                          .is_write_(QKV_is_write_out_31), .select_(QKV_selcet_out_31),
                          .calc_result_0(QKV_calc_result_31_0), .calc_result_1(QKV_calc_result_31_1), .calc_result_2(QKV_calc_result_31_2), .calc_result_3(QKV_calc_result_31_3), .calc_result_4(QKV_calc_result_31_4), .calc_result_5(QKV_calc_result_31_5), .calc_result_6(QKV_calc_result_31_6), .calc_result_7(QKV_calc_result_31_7), .calc_result_8(QKV_calc_result_31_8), .calc_result_9(QKV_calc_result_31_9), .calc_result_10(QKV_calc_result_31_10), .calc_result_11(QKV_calc_result_31_11), .calc_result_12(QKV_calc_result_31_12), .calc_result_13(QKV_calc_result_31_13), .calc_result_14(QKV_calc_result_31_14), .calc_result_15(QKV_calc_result_31_15)
);

dimc_macro i_dimc_macro_32(.input_addr(QKT_addr_out_0),
                          .input_weight_0(QKT_weight_out_0_0), .input_weight_1(QKT_weight_out_0_1), .input_weight_2(QKT_weight_out_0_2), .input_weight_3(QKT_weight_out_0_3), .input_weight_4(QKT_weight_out_0_4), .input_weight_5(QKT_weight_out_0_5), .input_weight_6(QKT_weight_out_0_6), .input_weight_7(QKT_weight_out_0_7), .input_weight_8(QKT_weight_out_0_8), .input_weight_9(QKT_weight_out_0_9), .input_weight_10(QKT_weight_out_0_10), .input_weight_11(QKT_weight_out_0_11), .input_weight_12(QKT_weight_out_0_12), .input_weight_13(QKT_weight_out_0_13), .input_weight_14(QKT_weight_out_0_14), .input_weight_15(QKT_weight_out_0_15),
                          .input_data_0(QKT_data_out_0_0), .input_data_1(QKT_data_out_0_1), .input_data_2(QKT_data_out_0_2), .input_data_3(QKT_data_out_0_3), .input_data_4(QKT_data_out_0_4), .input_data_5(QKT_data_out_0_5), .input_data_6(QKT_data_out_0_6), .input_data_7(QKT_data_out_0_7), .input_data_8(QKT_data_out_0_8), .input_data_9(QKT_data_out_0_9), .input_data_10(QKT_data_out_0_10), .input_data_11(QKT_data_out_0_11), .input_data_12(QKT_data_out_0_12), .input_data_13(QKT_data_out_0_13), .input_data_14(QKT_data_out_0_14), .input_data_15(QKT_data_out_0_15),
                          .is_write_(QKT_is_write_out_0), .select_(QKT_selcet_out_0),
                          .calc_result_0(QKT_calc_result_0_0), .calc_result_1(QKT_calc_result_0_1), .calc_result_2(QKT_calc_result_0_2), .calc_result_3(QKT_calc_result_0_3), .calc_result_4(QKT_calc_result_0_4), .calc_result_5(QKT_calc_result_0_5), .calc_result_6(QKT_calc_result_0_6), .calc_result_7(QKT_calc_result_0_7), .calc_result_8(QKT_calc_result_0_8), .calc_result_9(QKT_calc_result_0_9), .calc_result_10(QKT_calc_result_0_10), .calc_result_11(QKT_calc_result_0_11), .calc_result_12(QKT_calc_result_0_12), .calc_result_13(QKT_calc_result_0_13), .calc_result_14(QKT_calc_result_0_14), .calc_result_15(QKT_calc_result_0_15)
);

dimc_macro i_dimc_macro_33(.input_addr(QKT_addr_out_1),
                          .input_weight_0(QKT_weight_out_1_0), .input_weight_1(QKT_weight_out_1_1), .input_weight_2(QKT_weight_out_1_2), .input_weight_3(QKT_weight_out_1_3), .input_weight_4(QKT_weight_out_1_4), .input_weight_5(QKT_weight_out_1_5), .input_weight_6(QKT_weight_out_1_6), .input_weight_7(QKT_weight_out_1_7), .input_weight_8(QKT_weight_out_1_8), .input_weight_9(QKT_weight_out_1_9), .input_weight_10(QKT_weight_out_1_10), .input_weight_11(QKT_weight_out_1_11), .input_weight_12(QKT_weight_out_1_12), .input_weight_13(QKT_weight_out_1_13), .input_weight_14(QKT_weight_out_1_14), .input_weight_15(QKT_weight_out_1_15),
                          .input_data_0(QKT_data_out_1_0), .input_data_1(QKT_data_out_1_1), .input_data_2(QKT_data_out_1_2), .input_data_3(QKT_data_out_1_3), .input_data_4(QKT_data_out_1_4), .input_data_5(QKT_data_out_1_5), .input_data_6(QKT_data_out_1_6), .input_data_7(QKT_data_out_1_7), .input_data_8(QKT_data_out_1_8), .input_data_9(QKT_data_out_1_9), .input_data_10(QKT_data_out_1_10), .input_data_11(QKT_data_out_1_11), .input_data_12(QKT_data_out_1_12), .input_data_13(QKT_data_out_1_13), .input_data_14(QKT_data_out_1_14), .input_data_15(QKT_data_out_1_15),
                          .is_write_(QKT_is_write_out_1), .select_(QKT_selcet_out_1),
                          .calc_result_0(QKT_calc_result_1_0),

);

dimc_macro i_dimc_macro_34(.input_addr(QKT_addr_out_2),
                          .input_weight_0(QKT_weight_out_2_0), .input_weight_1(QKT_weight_out_2_1), .input_weight_2(QKT_weight_out_2_2), .input_weight_3(QKT_weight_out_2_3), .input_weight_4(QKT_weight_out_2_4), .input_weight_5(QKT_weight_out_2_5), .input_weight_6(QKT_weight_out_2_6), .input_weight_7(QKT_weight_out_2_7), .input_weight_8(QKT_weight_out_2_8), .input_weight_9(QKT_weight_out_2_9), .input_weight_10(QKT_weight_out_2_10), .input_weight_11(QKT_weight_out_2_11), .input_weight_12(QKT_weight_out_2_12), .input_weight_13(QKT_weight_out_2_13), .input_weight_14(QKT_weight_out_2_14), .input_weight_15(QKT_weight_out_2_15),
                          .input_data_0(QKT_data_out_2_0), .input_data_1(QKT_data_out_2_1), .input_data_2(QKT_data_out_2_2), .input_data_3(QKT_data_out_2_3), .input_data_4(QKT_data_out_2_4), .input_data_5(QKT_data_out_2_5), .input_data_6(QKT_data_out_2_6), .input_data_7(QKT_data_out_2_7), .input_data_8(QKT_data_out_2_8), .input_data_9(QKT_data_out_2_9), .input_data_10(QKT_data_out_2_10), .input_data_11(QKT_data_out_2_11), .input_data_12(QKT_data_out_2_12), .input_data_13(QKT_data_out_2_13), .input_data_14(QKT_data_out_2_14), .input_data_15(QKT_data_out_2_15),
                          .is_write_(QKT_is_write_out_2), .select_(QKT_selcet_out_2),
                          .calc_result_0(QKT_calc_result_2_0),

);

dimc_macro i_dimc_macro_35(.input_addr(QKT_addr_out_3),
                          .input_weight_0(QKT_weight_out_3_0), .input_weight_1(QKT_weight_out_3_1), .input_weight_2(QKT_weight_out_3_2), .input_weight_3(QKT_weight_out_3_3), .input_weight_4(QKT_weight_out_3_4), .input_weight_5(QKT_weight_out_3_5), .input_weight_6(QKT_weight_out_3_6), .input_weight_7(QKT_weight_out_3_7), .input_weight_8(QKT_weight_out_3_8), .input_weight_9(QKT_weight_out_3_9), .input_weight_10(QKT_weight_out_3_10), .input_weight_11(QKT_weight_out_3_11), .input_weight_12(QKT_weight_out_3_12), .input_weight_13(QKT_weight_out_3_13), .input_weight_14(QKT_weight_out_3_14), .input_weight_15(QKT_weight_out_3_15),
                          .input_data_0(QKT_data_out_3_0), .input_data_1(QKT_data_out_3_1), .input_data_2(QKT_data_out_3_2), .input_data_3(QKT_data_out_3_3), .input_data_4(QKT_data_out_3_4), .input_data_5(QKT_data_out_3_5), .input_data_6(QKT_data_out_3_6), .input_data_7(QKT_data_out_3_7), .input_data_8(QKT_data_out_3_8), .input_data_9(QKT_data_out_3_9), .input_data_10(QKT_data_out_3_10), .input_data_11(QKT_data_out_3_11), .input_data_12(QKT_data_out_3_12), .input_data_13(QKT_data_out_3_13), .input_data_14(QKT_data_out_3_14), .input_data_15(QKT_data_out_3_15),
                          .is_write_(QKT_is_write_out_3), .select_(QKT_selcet_out_3),
                          .calc_result_0(QKT_calc_result_3_0),

);

endmodule
